//Verilog HDL for "Lib6710_08", "TIELO" "functional"


module TIELO ( Y );

  output Y;
   assign Y = 0;
   
endmodule
