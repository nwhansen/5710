/home/nathan/5710/libfiles/11-17/Lib6710_08.lef