//Verilog HDL for "Lib6710_08", "AOI22X1" "functional"


module AOI22X1 ( );

endmodule
