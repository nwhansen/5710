/home/nathan/5710/libfiles/current/Lib6710_08.lef