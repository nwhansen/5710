// Global nets module 

`celldefine
module cds_globals;



endmodule
`endcelldefine
