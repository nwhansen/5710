//Verilog HDL for "lab5", "tiehi" "behavioral"


module TIEHI(Y);
  output Y;
  assign Y = 1;
endmodule
