###########################
# 
# This is the TechHeader.lef file that contains the 
# technology information for the AMI C5N 0.5 micron 
# CMOS technology (SCN3M_SUBM when using MOSIS)
# 
# Erik Brunvand
###########################

VERSION 5.6 ;

BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
  LIBRARY minWidth REAL 1.5 ;
  LIBRARY PadType STRING "Perimeter" ;
  LIBRARY technology STRING "UofU_AMI_C5N" ;
  LIBRARY model STRING "ami06" ;
  LIBRARY gridResolution REAL 0.15 ;
  LIBRARY minLength REAL 0.6 ;
  LAYER sheetResistance INTEGER ;
END PROPERTYDEFINITIONS

UNITS
  DATABASE MICRONS 1000 ;
END UNITS
MANUFACTURINGGRID 0.15 ;

LAYER poly
  TYPE  MASTERSLICE ;
END poly

LAYER cc
  TYPE  CUT ;
  SPACING       0.9 ;
END cc

LAYER metal1
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3 3 ;
  WIDTH 0.9 ;
  SPACING 0.9 ;
  OFFSET 1.5 ;
  THICKNESS 0.64 ;
  HEIGHT 0.38 ;
  RESISTANCE RPERSQ 0.09 ;
  CAPACITANCE CPERSQDIST 3.2e-05 ;
  EDGECAPACITANCE 7.5e-05 ;
END metal1

LAYER via
  TYPE CUT ;
  SPACING 0.9 ;
END via

LAYER metal2
  TYPE ROUTING ;
  DIRECTION VERTICAL ;
  PITCH 2.4 2.4 ;
  WIDTH 0.9 ;
  SPACING 0.9 ;
  OFFSET        1.2 ;
  THICKNESS 0.57 ;
  HEIGHT 1.62 ;
  RESISTANCE RPERSQ 0.09 ;
  CAPACITANCE CPERSQDIST 1.6e-05 ;
  EDGECAPACITANCE 6.0e-05 ;
END metal2

LAYER via2
  TYPE CUT ;
  SPACING 0.9 ;
END via2

LAYER metal3
  TYPE ROUTING ;
  DIRECTION HORIZONTAL ;
  PITCH 3 3 ;
  WIDTH 1.5 ;
  SPACING 0.9 ;
  OFFSET        1.5 ;
  THICKNESS 0.77 ;
  HEIGHT 2.52 ;
  RESISTANCE RPERSQ 0.05 ;
  CAPACITANCE CPERSQDIST 1e-05 ;
  EDGECAPACITANCE 4.0e-05 ;
END metal3

LAYER OVERLAP
  TYPE OVERLAP ;
END OVERLAP

VIA M2_M1_via DEFAULT
  LAYER metal1 ;
    RECT -0.6 -0.6 0.6 0.6 ;
  LAYER via ;
    RECT -0.3 -0.3 0.3 0.3 ;
  LAYER metal2 ;
    RECT -0.6 -0.6 0.6 0.6 ;
END M2_M1_via

VIA M3_M2_via DEFAULT
  LAYER metal2 ;
    RECT -0.6 -0.6 0.6 0.6 ;
  LAYER via2 ;
    RECT -0.3 -0.3 0.3 0.3 ;
  LAYER metal3 ;
    RECT -0.9 -0.9 0.9 0.9 ;
END M3_M2_via

VIARULE M3_M2 GENERATE
  LAYER metal2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER metal3 ;
    ENCLOSURE 0.6 0.6 ;
  LAYER via2 ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.5 BY 1.5 ;
END M3_M2

VIARULE M2_M1 GENERATE
  LAYER metal1 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER metal2 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER via ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.5 BY 1.5 ;
END M2_M1

VIARULE viagen21 GENERATE
  LAYER metal1 ;
    WIDTH 1.2 TO 120 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER metal2 ;
    WIDTH 1.2 TO 120 ;
    ENCLOSURE 0.3 0.3 ;
  LAYER via ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 1.5 BY 1.5 ;
END viagen21

VIARULE viagen32 GENERATE
  LAYER metal2 ;
    WIDTH 1.2 TO 120 ;
    ENCLOSURE 0.6 0.6 ;
  LAYER metal3 ;
    WIDTH 1.8 TO 180 ;
    ENCLOSURE 0.6 0.6 ;
  LAYER via2 ;
    RECT -0.3 -0.3 0.3 0.3 ;
    SPACING 2.1 BY 2.1 ;
END viagen32

#SPACING
#  SAMENET metal1 metal1 0.9 ;
#  SAMENET metal2 metal2 0.9 ;
#  SAMENET metal3 metal3 0.9 ;
#END SPACING

SPACING
  SAMENET metal1  metal1        0.900  STACK ;
  SAMENET metal2  metal2        0.900  STACK ;
  SAMENET metal3  metal3        0.900 ;
  SAMENET cc  via       0.000  STACK ;
  SAMENET via  via      0.900 ;
  SAMENET via  via2     0.000  STACK ;
  SAMENET via2  via2    0.900 ;
END SPACING

SITE corner
  CLASS PAD ;
  SYMMETRY Y R90 ;
  SIZE 300 BY 300 ;
END corner

SITE IO
  CLASS PAD ;
  SYMMETRY Y ;
  SIZE 90 BY 300 ;
END IO

SITE  dbl_core
    CLASS       CORE ;
    SYMMETRY    Y ;
    SIZE        2.400 BY 54.000 ;
END  dbl_core

SITE core
  CLASS CORE ;
  SYMMETRY Y ;
  SIZE 2.4 BY 27 ;
END core

MACRO XOR2X1
    CLASS CORE ;
    FOREIGN XOR2X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.20 3.90 13.80 ;
        LAYER metal2 ;
        RECT  3.00 12.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 12.90 4.20 14.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 18.00 6.30 18.60 ;
        LAYER metal2 ;
        RECT  5.40 6.60 6.60 18.90 ;
        LAYER metal1 ;
        RECT  5.40 5.10 8.40 6.30 ;
        RECT  7.20 2.10 8.40 6.30 ;
        RECT  5.40 5.10 6.60 7.80 ;
        RECT  6.90 17.70 8.10 24.90 ;
        RECT  5.40 17.70 8.10 18.90 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  12.90 12.90 13.50 13.50 ;
        LAYER metal2 ;
        RECT  12.60 12.60 13.80 14.10 ;
        LAYER metal1 ;
        RECT  12.60 12.60 13.80 13.80 ;
        RECT  7.80 12.60 13.80 13.50 ;
        RECT  7.80 12.30 9.00 13.50 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 18.00 1.20 ;
        RECT  11.10 -1.20 12.30 7.50 ;
        RECT  3.00 -1.20 4.20 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 18.00 28.20 ;
        RECT  11.10 16.50 12.30 28.20 ;
        RECT  3.00 16.50 4.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 16.80 3.90 17.40 ;
        RECT  3.30 13.20 3.90 13.80 ;
        RECT  3.30 6.60 3.90 7.20 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  6.60 15.00 7.20 15.60 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 24.00 7.80 24.60 ;
        RECT  7.20 22.50 7.80 23.10 ;
        RECT  7.20 21.00 7.80 21.60 ;
        RECT  7.20 19.50 7.80 20.10 ;
        RECT  7.20 18.00 7.80 18.60 ;
        RECT  7.50 5.40 8.10 6.00 ;
        RECT  7.50 3.90 8.10 4.50 ;
        RECT  7.50 2.40 8.10 3.00 ;
        RECT  8.10 12.60 8.70 13.20 ;
        RECT  8.10 8.70 8.70 9.30 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.50 10.80 11.10 11.40 ;
        RECT  11.40 24.30 12.00 24.90 ;
        RECT  11.40 22.80 12.00 23.40 ;
        RECT  11.40 21.30 12.00 21.90 ;
        RECT  11.40 19.80 12.00 20.40 ;
        RECT  11.40 18.30 12.00 18.90 ;
        RECT  11.40 16.80 12.00 17.40 ;
        RECT  11.40 6.60 12.00 7.20 ;
        RECT  11.40 5.10 12.00 5.70 ;
        RECT  11.40 3.60 12.00 4.20 ;
        RECT  11.40 2.10 12.00 2.70 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.90 12.90 13.50 13.50 ;
        RECT  13.80 24.00 14.40 24.60 ;
        RECT  13.80 22.50 14.40 23.10 ;
        RECT  13.80 21.00 14.40 21.60 ;
        RECT  13.80 19.50 14.40 20.10 ;
        RECT  13.80 3.90 14.40 4.50 ;
        RECT  13.80 2.40 14.40 3.00 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        LAYER metal1 ;
        RECT  0.60 10.50 11.40 11.40 ;
        RECT  10.20 10.50 11.40 11.70 ;
        RECT  0.60 2.10 1.80 24.90 ;
        RECT  13.50 2.10 15.90 4.80 ;
        RECT  7.80 8.40 15.90 9.60 ;
        RECT  6.30 14.70 15.90 15.60 ;
        RECT  6.30 14.70 7.50 15.90 ;
        RECT  14.70 2.10 15.90 24.90 ;
        RECT  13.50 19.20 15.90 24.90 ;
    END
END XOR2X1

MACRO XNOR2X1
    CLASS CORE ;
    FOREIGN XNOR2X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.20 3.90 13.80 ;
        LAYER metal2 ;
        RECT  3.00 12.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 12.90 4.20 14.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 18.00 6.30 18.60 ;
        LAYER metal2 ;
        RECT  5.40 6.60 6.60 18.90 ;
        LAYER metal1 ;
        RECT  5.40 5.10 8.40 6.30 ;
        RECT  7.20 2.10 8.40 6.30 ;
        RECT  5.40 5.10 6.60 7.80 ;
        RECT  6.90 17.70 8.10 24.90 ;
        RECT  5.40 17.70 8.10 18.90 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  12.90 9.90 13.50 10.50 ;
        LAYER metal2 ;
        RECT  12.60 9.60 13.80 11.10 ;
        LAYER metal1 ;
        RECT  12.60 8.40 13.80 10.80 ;
        RECT  7.80 8.40 13.80 9.60 ;
        END
    END B
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 18.00 1.20 ;
        RECT  11.10 -1.20 12.30 7.50 ;
        RECT  3.00 -1.20 4.20 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 18.00 28.20 ;
        RECT  11.10 16.50 12.30 28.20 ;
        RECT  3.00 16.50 4.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 16.80 3.90 17.40 ;
        RECT  3.30 13.20 3.90 13.80 ;
        RECT  3.30 6.60 3.90 7.20 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  6.60 15.00 7.20 15.60 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 24.00 7.80 24.60 ;
        RECT  7.20 22.50 7.80 23.10 ;
        RECT  7.20 21.00 7.80 21.60 ;
        RECT  7.20 19.50 7.80 20.10 ;
        RECT  7.20 18.00 7.80 18.60 ;
        RECT  7.50 5.40 8.10 6.00 ;
        RECT  7.50 3.90 8.10 4.50 ;
        RECT  7.50 2.40 8.10 3.00 ;
        RECT  8.10 12.60 8.70 13.20 ;
        RECT  8.10 8.70 8.70 9.30 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.50 10.80 11.10 11.40 ;
        RECT  11.40 24.30 12.00 24.90 ;
        RECT  11.40 22.80 12.00 23.40 ;
        RECT  11.40 21.30 12.00 21.90 ;
        RECT  11.40 19.80 12.00 20.40 ;
        RECT  11.40 18.30 12.00 18.90 ;
        RECT  11.40 16.80 12.00 17.40 ;
        RECT  11.40 6.60 12.00 7.20 ;
        RECT  11.40 5.10 12.00 5.70 ;
        RECT  11.40 3.60 12.00 4.20 ;
        RECT  11.40 2.10 12.00 2.70 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.75 14.70 13.35 15.30 ;
        RECT  12.90 9.90 13.50 10.50 ;
        RECT  13.80 24.00 14.40 24.60 ;
        RECT  13.80 22.50 14.40 23.10 ;
        RECT  13.80 21.00 14.40 21.60 ;
        RECT  13.80 19.50 14.40 20.10 ;
        RECT  13.80 3.90 14.40 4.50 ;
        RECT  13.80 2.40 14.40 3.00 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        LAYER metal1 ;
        RECT  0.60 10.50 11.40 11.40 ;
        RECT  10.20 10.50 11.40 11.70 ;
        RECT  0.60 2.10 1.80 24.90 ;
        RECT  12.45 14.40 13.65 15.60 ;
        RECT  6.30 14.70 13.65 15.60 ;
        RECT  6.30 14.70 7.50 15.90 ;
        RECT  13.50 2.10 15.90 4.80 ;
        RECT  7.80 12.30 9.00 13.50 ;
        RECT  7.80 12.60 15.90 13.50 ;
        RECT  14.70 2.10 15.90 24.90 ;
        RECT  13.50 19.20 15.90 24.90 ;
    END
END XNOR2X1

MACRO TIELO
    CLASS CORE ;
    FOREIGN TIELO 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 5.10 ;
        LAYER metal1 ;
        RECT  3.00 2.10 4.20 5.10 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 6.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 6.00 1.20 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 17.70 3.90 18.30 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        LAYER metal1 ;
        RECT  3.00 17.40 4.20 24.90 ;
    END
END TIELO

MACRO TIEHI
    CLASS CORE ;
    FOREIGN TIEHI 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        LAYER metal2 ;
        RECT  3.00 19.20 4.20 24.90 ;
        LAYER metal1 ;
        RECT  3.00 19.20 4.20 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 6.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 6.00 1.20 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 5.70 3.90 6.30 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        LAYER metal1 ;
        RECT  3.00 2.10 4.20 6.60 ;
    END
END TIEHI

MACRO OAI22X1
    CLASS CORE ;
    FOREIGN OAI22X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 18.90 ;
        LAYER metal1 ;
        RECT  5.40 13.20 6.60 24.90 ;
        RECT  3.00 13.20 6.60 18.90 ;
        RECT  3.00 2.10 4.20 4.80 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  7.20 7.80 7.80 8.40 ;
        LAYER metal2 ;
        RECT  6.90 7.50 9.00 8.70 ;
        RECT  7.80 6.90 9.00 8.70 ;
        LAYER metal1 ;
        RECT  6.90 7.50 8.10 8.70 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  10.50 10.20 11.10 10.80 ;
        LAYER metal2 ;
        RECT  10.20 3.90 11.40 11.10 ;
        LAYER metal1 ;
        RECT  10.20 9.90 11.40 11.10 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 10.20 6.30 10.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  4.50 9.90 6.60 11.10 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 12.00 1.50 12.60 ;
        LAYER metal2 ;
        RECT  0.60 11.70 1.80 14.10 ;
        LAYER metal1 ;
        RECT  0.60 11.70 1.80 12.90 ;
        END
    END D
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 13.20 28.20 ;
        RECT  9.45 13.50 10.65 28.20 ;
        RECT  0.90 15.00 2.10 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 13.20 1.20 ;
        RECT  7.80 -1.20 9.00 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 12.00 1.50 12.60 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  1.20 24.30 1.80 24.90 ;
        RECT  1.20 22.80 1.80 23.40 ;
        RECT  1.20 21.30 1.80 21.90 ;
        RECT  1.20 19.80 1.80 20.40 ;
        RECT  1.20 18.30 1.80 18.90 ;
        RECT  1.20 16.80 1.80 17.40 ;
        RECT  1.20 15.30 1.80 15.90 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 10.20 5.40 10.80 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 18.00 6.30 18.60 ;
        RECT  5.70 16.50 6.30 17.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 13.50 6.30 14.10 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 7.80 7.80 8.40 ;
        RECT  8.10 3.60 8.70 4.20 ;
        RECT  8.10 2.10 8.70 2.70 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  9.75 24.30 10.35 24.90 ;
        RECT  9.75 22.80 10.35 23.40 ;
        RECT  9.75 21.30 10.35 21.90 ;
        RECT  9.75 19.80 10.35 20.40 ;
        RECT  9.75 18.30 10.35 18.90 ;
        RECT  9.75 16.80 10.35 17.40 ;
        RECT  9.75 15.30 10.35 15.90 ;
        RECT  9.75 13.80 10.35 14.40 ;
        RECT  10.50 10.20 11.10 10.80 ;
        RECT  10.50 3.90 11.10 4.50 ;
        RECT  10.50 2.40 11.10 3.00 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        LAYER metal1 ;
        RECT  0.60 2.10 1.80 6.60 ;
        RECT  5.40 2.10 6.60 6.60 ;
        RECT  10.20 2.10 11.40 6.60 ;
        RECT  0.60 5.70 11.40 6.60 ;
    END
END OAI22X1

MACRO OAI21X1
    CLASS CORE ;
    FOREIGN OAI21X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 10.20 6.30 10.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  3.90 9.90 6.60 11.10 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 6.90 9.00 11.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 9.00 11.10 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 16.20 1.50 16.80 ;
        LAYER metal2 ;
        RECT  0.60 15.90 1.80 17.10 ;
        LAYER metal1 ;
        RECT  0.60 15.90 1.80 17.10 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        LAYER metal2 ;
        RECT  3.00 13.20 4.20 18.90 ;
        LAYER metal1 ;
        RECT  3.00 12.00 4.20 24.90 ;
        RECT  0.60 12.00 4.20 13.20 ;
        RECT  0.60 2.10 1.80 13.20 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 10.80 28.20 ;
        RECT  6.90 13.50 8.10 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 10.80 1.20 ;
        RECT  5.40 -1.20 6.60 6.00 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 16.20 1.50 16.80 ;
        RECT  0.90 6.90 1.50 7.50 ;
        RECT  0.90 5.40 1.50 6.00 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.20 10.20 4.80 10.80 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 5.10 6.30 5.70 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 24.30 7.80 24.90 ;
        RECT  7.20 22.80 7.80 23.40 ;
        RECT  7.20 21.30 7.80 21.90 ;
        RECT  7.20 19.80 7.80 20.40 ;
        RECT  7.20 18.30 7.80 18.90 ;
        RECT  7.20 16.80 7.80 17.40 ;
        RECT  7.20 15.30 7.80 15.90 ;
        RECT  7.20 13.80 7.80 14.40 ;
        RECT  8.10 10.20 8.70 10.80 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        LAYER metal1 ;
        RECT  3.00 2.10 4.20 8.10 ;
        RECT  7.80 2.10 9.00 8.10 ;
        RECT  3.00 6.90 9.00 8.10 ;
    END
END OAI21X1

MACRO NOR3X1
    CLASS CORE ;
    FOREIGN NOR3X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  15.30 10.20 15.90 10.80 ;
        LAYER metal2 ;
        RECT  15.00 9.90 16.20 14.40 ;
        LAYER metal1 ;
        RECT  15.00 9.90 16.20 11.10 ;
        END
    END C
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 11.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 9.00 11.10 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 7.20 3.90 7.80 ;
        LAYER metal2 ;
        RECT  3.00 6.90 4.20 8.10 ;
        LAYER metal1 ;
        RECT  3.00 6.90 4.20 8.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  17.70 22.50 18.30 23.10 ;
        LAYER metal2 ;
        RECT  17.40 22.20 18.60 23.40 ;
        LAYER metal1 ;
        RECT  17.40 13.50 18.60 23.40 ;
        RECT  12.60 13.50 18.60 14.40 ;
        RECT  8.70 5.55 14.70 6.45 ;
        RECT  13.50 2.10 14.70 6.45 ;
        RECT  12.60 5.55 13.80 21.90 ;
        RECT  8.70 2.10 9.90 6.45 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 20.40 28.20 ;
        RECT  3.00 16.20 4.20 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 20.40 1.20 ;
        RECT  11.10 -1.20 12.30 4.50 ;
        RECT  6.30 -1.20 7.50 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 18.00 1.50 18.60 ;
        RECT  0.90 16.50 1.50 17.10 ;
        RECT  0.90 15.00 1.50 15.60 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 16.80 3.90 17.40 ;
        RECT  3.30 7.20 3.90 7.80 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 18.00 6.30 18.60 ;
        RECT  5.70 16.50 6.30 17.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  6.60 3.60 7.20 4.20 ;
        RECT  6.60 2.10 7.20 2.70 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 10.20 8.70 10.80 ;
        RECT  9.00 3.90 9.60 4.50 ;
        RECT  9.00 2.40 9.60 3.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.50 21.00 11.10 21.60 ;
        RECT  10.50 19.50 11.10 20.10 ;
        RECT  10.50 18.00 11.10 18.60 ;
        RECT  10.50 16.50 11.10 17.10 ;
        RECT  10.50 15.00 11.10 15.60 ;
        RECT  11.40 3.60 12.00 4.20 ;
        RECT  11.40 2.10 12.00 2.70 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.90 21.00 13.50 21.60 ;
        RECT  12.90 19.50 13.50 20.10 ;
        RECT  12.90 18.00 13.50 18.60 ;
        RECT  12.90 16.50 13.50 17.10 ;
        RECT  12.90 15.00 13.50 15.60 ;
        RECT  13.80 3.90 14.40 4.50 ;
        RECT  13.80 2.40 14.40 3.00 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.30 22.50 15.90 23.10 ;
        RECT  15.30 21.00 15.90 21.60 ;
        RECT  15.30 19.50 15.90 20.10 ;
        RECT  15.30 18.00 15.90 18.60 ;
        RECT  15.30 16.50 15.90 17.10 ;
        RECT  15.30 10.20 15.90 10.80 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 22.50 18.30 23.10 ;
        RECT  17.70 21.00 18.30 21.60 ;
        RECT  17.70 19.50 18.30 20.10 ;
        RECT  17.70 18.00 18.30 18.60 ;
        RECT  17.70 16.50 18.30 17.10 ;
        RECT  17.70 15.00 18.30 15.60 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        LAYER metal1 ;
        RECT  0.60 13.50 11.40 14.40 ;
        RECT  10.20 13.50 11.40 21.90 ;
        RECT  0.60 13.50 1.80 23.40 ;
        RECT  5.40 13.50 6.60 23.40 ;
        RECT  7.80 16.20 9.00 24.90 ;
        RECT  15.00 16.20 16.20 24.90 ;
        RECT  7.80 24.00 16.20 24.90 ;
    END
END NOR3X1

MACRO NOR2X2
    CLASS CORE ;
    FOREIGN NOR2X2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 12.00 3.90 12.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 14.40 ;
        LAYER metal1 ;
        RECT  4.50 13.20 5.70 23.40 ;
        RECT  3.00 13.20 5.70 14.40 ;
        RECT  3.00 11.70 4.20 14.40 ;
        RECT  3.00 2.10 4.20 7.80 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 9.00 6.30 9.60 ;
        LAYER metal2 ;
        RECT  5.40 8.70 6.60 14.10 ;
        LAYER metal1 ;
        RECT  5.40 8.70 6.60 9.90 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 13.20 28.20 ;
        RECT  8.40 13.80 9.60 28.20 ;
        RECT  0.60 13.80 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 13.20 1.20 ;
        RECT  5.40 -1.20 6.60 7.50 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 23.10 1.50 23.70 ;
        RECT  0.90 21.60 1.50 22.20 ;
        RECT  0.90 20.10 1.50 20.70 ;
        RECT  0.90 18.60 1.50 19.20 ;
        RECT  0.90 17.10 1.50 17.70 ;
        RECT  0.90 15.60 1.50 16.20 ;
        RECT  0.90 14.10 1.50 14.70 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 22.50 5.40 23.10 ;
        RECT  4.80 21.00 5.40 21.60 ;
        RECT  4.80 19.50 5.40 20.10 ;
        RECT  4.80 18.00 5.40 18.60 ;
        RECT  4.80 16.50 5.40 17.10 ;
        RECT  4.80 15.00 5.40 15.60 ;
        RECT  4.80 13.50 5.40 14.10 ;
        RECT  5.70 9.00 6.30 9.60 ;
        RECT  5.70 6.60 6.30 7.20 ;
        RECT  5.70 5.10 6.30 5.70 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.70 23.10 9.30 23.70 ;
        RECT  8.70 21.60 9.30 22.20 ;
        RECT  8.70 20.10 9.30 20.70 ;
        RECT  8.70 18.60 9.30 19.20 ;
        RECT  8.70 17.10 9.30 17.70 ;
        RECT  8.70 15.60 9.30 16.20 ;
        RECT  8.70 14.10 9.30 14.70 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
    END
END NOR2X2

MACRO NOR2X1
    CLASS CORE ;
    FOREIGN NOR2X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 12.00 3.90 12.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 14.40 ;
        LAYER metal1 ;
        RECT  4.50 13.20 5.70 24.90 ;
        RECT  3.00 13.20 5.70 14.40 ;
        RECT  3.00 11.70 4.20 14.40 ;
        RECT  3.00 2.10 4.20 4.80 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 7.20 1.50 7.80 ;
        LAYER metal2 ;
        RECT  0.60 6.90 1.80 8.10 ;
        LAYER metal1 ;
        RECT  0.60 6.90 1.80 8.10 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 10.20 6.30 10.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  5.40 9.90 6.60 11.10 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 8.40 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 8.40 1.20 ;
        RECT  5.40 -1.20 6.60 4.50 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  0.90 7.20 1.50 7.80 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 24.00 5.40 24.60 ;
        RECT  4.80 22.50 5.40 23.10 ;
        RECT  4.80 21.00 5.40 21.60 ;
        RECT  4.80 19.50 5.40 20.10 ;
        RECT  4.80 18.00 5.40 18.60 ;
        RECT  4.80 16.50 5.40 17.10 ;
        RECT  4.80 15.00 5.40 15.60 ;
        RECT  4.80 13.50 5.40 14.10 ;
        RECT  5.70 10.20 6.30 10.80 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
    END
END NOR2X1

MACRO NAND3X1
    CLASS CORE ;
    FOREIGN NAND3X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 15.60 3.90 16.20 ;
        LAYER metal2 ;
        RECT  3.00 15.30 4.20 20.10 ;
        LAYER metal1 ;
        RECT  3.00 15.30 4.20 16.50 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 13.20 6.30 13.80 ;
        LAYER metal2 ;
        RECT  5.40 12.90 6.60 14.10 ;
        LAYER metal1 ;
        RECT  5.40 12.90 6.60 14.10 ;
        END
    END B
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 11.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 10.50 11.10 ;
        RECT  9.30 2.10 10.50 11.10 ;
        RECT  7.80 9.90 9.00 24.90 ;
        RECT  3.00 17.40 9.00 18.60 ;
        RECT  3.00 17.40 4.20 24.90 ;
        END
    END Y
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  10.50 16.20 11.10 16.80 ;
        LAYER metal2 ;
        RECT  10.20 15.90 11.40 17.10 ;
        LAYER metal1 ;
        RECT  10.20 15.90 11.40 17.10 ;
        END
    END C
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 15.60 28.20 ;
        RECT  10.20 19.50 11.40 28.20 ;
        RECT  5.40 19.50 6.60 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 15.60 1.20 ;
        RECT  3.90 -1.20 5.10 10.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 15.60 3.90 16.20 ;
        RECT  4.20 9.60 4.80 10.20 ;
        RECT  4.20 8.10 4.80 8.70 ;
        RECT  4.20 6.60 4.80 7.20 ;
        RECT  4.20 5.10 4.80 5.70 ;
        RECT  4.20 3.60 4.80 4.20 ;
        RECT  4.20 2.10 4.80 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 13.20 6.30 13.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  9.60 9.90 10.20 10.50 ;
        RECT  9.60 8.40 10.20 9.00 ;
        RECT  9.60 6.90 10.20 7.50 ;
        RECT  9.60 5.40 10.20 6.00 ;
        RECT  9.60 3.90 10.20 4.50 ;
        RECT  9.60 2.40 10.20 3.00 ;
        RECT  10.50 24.30 11.10 24.90 ;
        RECT  10.50 22.80 11.10 23.40 ;
        RECT  10.50 21.30 11.10 21.90 ;
        RECT  10.50 19.80 11.10 20.40 ;
        RECT  10.50 16.20 11.10 16.80 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
    END
END NAND3X1

MACRO NAND2X2
    CLASS CORE ;
    FOREIGN NAND2X2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 14.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        LAYER metal2 ;
        RECT  3.00 3.60 4.20 24.90 ;
        LAYER metal1 ;
        RECT  4.50 3.00 5.70 8.70 ;
        RECT  3.00 3.60 5.70 7.80 ;
        RECT  3.00 13.20 4.20 24.90 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 10.20 6.30 10.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  4.20 9.90 6.60 11.10 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 13.20 28.20 ;
        RECT  5.40 13.50 6.60 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 13.20 1.20 ;
        RECT  8.40 -1.20 9.60 8.70 ;
        RECT  0.60 -1.20 1.80 8.70 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 7.80 1.50 8.40 ;
        RECT  0.90 6.30 1.50 6.90 ;
        RECT  0.90 4.80 1.50 5.40 ;
        RECT  0.90 3.30 1.50 3.90 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 10.20 5.10 10.80 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 7.80 5.40 8.40 ;
        RECT  4.80 6.30 5.40 6.90 ;
        RECT  4.80 4.80 5.40 5.40 ;
        RECT  4.80 3.30 5.40 3.90 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 18.30 6.30 18.90 ;
        RECT  5.70 16.80 6.30 17.40 ;
        RECT  5.70 15.30 6.30 15.90 ;
        RECT  5.70 13.80 6.30 14.40 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.70 7.80 9.30 8.40 ;
        RECT  8.70 6.30 9.30 6.90 ;
        RECT  8.70 4.80 9.30 5.40 ;
        RECT  8.70 3.30 9.30 3.90 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
    END
END NAND2X2

MACRO NAND2X1
    CLASS CORE ;
    FOREIGN NAND2X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 13.20 1.50 13.80 ;
        LAYER metal2 ;
        RECT  0.60 12.90 1.80 14.10 ;
        LAYER metal1 ;
        RECT  0.60 12.90 1.80 14.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 8.40 3.90 9.00 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        LAYER metal2 ;
        RECT  3.00 6.60 4.20 24.90 ;
        LAYER metal1 ;
        RECT  3.00 6.60 5.70 7.80 ;
        RECT  4.50 2.10 5.70 7.80 ;
        RECT  3.00 6.60 4.20 9.30 ;
        RECT  3.00 19.20 4.20 24.90 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 10.20 6.30 10.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  5.40 9.90 6.60 11.10 ;
        END
    END B
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 8.40 28.20 ;
        RECT  5.40 19.50 6.60 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 8.40 1.20 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 13.20 1.50 13.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 6.90 5.40 7.50 ;
        RECT  4.80 5.40 5.40 6.00 ;
        RECT  4.80 3.90 5.40 4.50 ;
        RECT  4.80 2.40 5.40 3.00 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 10.20 6.30 10.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
    END
END NAND2X1

MACRO MUX2X2
    CLASS CORE ;
    FOREIGN MUX2X2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 19.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 13.20 6.30 13.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 14.10 ;
        LAYER metal1 ;
        RECT  5.40 12.90 6.60 14.10 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  12.90 12.90 13.50 13.50 ;
        LAYER metal2 ;
        RECT  12.60 12.60 13.80 17.10 ;
        LAYER metal1 ;
        RECT  9.60 12.60 13.80 13.80 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.20 3.90 13.80 ;
        LAYER metal2 ;
        RECT  3.00 12.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 12.90 4.20 14.10 ;
        END
    END S
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  15.90 13.50 16.50 14.10 ;
        RECT  15.90 15.00 16.50 15.60 ;
        RECT  15.90 16.50 16.50 17.10 ;
        RECT  15.90 18.00 16.50 18.60 ;
        RECT  15.90 19.50 16.50 20.10 ;
        RECT  15.90 21.00 16.50 21.60 ;
        RECT  15.90 22.50 16.50 23.10 ;
        RECT  15.90 24.00 16.50 24.60 ;
        LAYER metal2 ;
        RECT  15.60 13.20 16.80 24.90 ;
        LAYER metal1 ;
        RECT  15.60 2.10 16.80 24.90 ;
        END
    END Y
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 20.40 1.20 ;
        RECT  12.60 -1.20 13.80 6.00 ;
        RECT  3.00 -1.20 5.70 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 20.40 28.20 ;
        RECT  12.60 18.00 13.80 28.20 ;
        RECT  3.00 18.00 5.70 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.00 10.80 3.60 11.40 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 13.20 3.90 13.80 ;
        RECT  3.30 6.60 3.90 7.20 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 24.30 5.40 24.90 ;
        RECT  4.80 22.80 5.40 23.40 ;
        RECT  4.80 21.30 5.40 21.90 ;
        RECT  4.80 19.80 5.40 20.40 ;
        RECT  4.80 18.30 5.40 18.90 ;
        RECT  4.80 6.60 5.40 7.20 ;
        RECT  4.80 5.10 5.40 5.70 ;
        RECT  4.80 3.60 5.40 4.20 ;
        RECT  4.80 2.10 5.40 2.70 ;
        RECT  5.40 8.70 6.00 9.30 ;
        RECT  5.70 13.20 6.30 13.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  9.00 24.00 9.60 24.60 ;
        RECT  9.00 22.50 9.60 23.10 ;
        RECT  9.00 21.00 9.60 21.60 ;
        RECT  9.00 19.50 9.60 20.10 ;
        RECT  9.00 18.00 9.60 18.60 ;
        RECT  9.00 6.90 9.60 7.50 ;
        RECT  9.00 5.40 9.60 6.00 ;
        RECT  9.00 3.90 9.60 4.50 ;
        RECT  9.00 2.40 9.60 3.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  9.90 12.90 10.50 13.50 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.30 15.00 12.90 15.60 ;
        RECT  12.30 10.80 12.90 11.40 ;
        RECT  12.90 24.30 13.50 24.90 ;
        RECT  12.90 22.80 13.50 23.40 ;
        RECT  12.90 21.30 13.50 21.90 ;
        RECT  12.90 19.80 13.50 20.40 ;
        RECT  12.90 18.30 13.50 18.90 ;
        RECT  12.90 5.10 13.50 5.70 ;
        RECT  12.90 3.60 13.50 4.20 ;
        RECT  12.90 2.10 13.50 2.70 ;
        RECT  13.80 8.40 14.40 9.00 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.90 24.00 16.50 24.60 ;
        RECT  15.90 22.50 16.50 23.10 ;
        RECT  15.90 21.00 16.50 21.60 ;
        RECT  15.90 19.50 16.50 20.10 ;
        RECT  15.90 18.00 16.50 18.60 ;
        RECT  15.90 16.50 16.50 17.10 ;
        RECT  15.90 15.00 16.50 15.60 ;
        RECT  15.90 13.50 16.50 14.10 ;
        RECT  15.90 6.90 16.50 7.50 ;
        RECT  15.90 5.40 16.50 6.00 ;
        RECT  15.90 3.90 16.50 4.50 ;
        RECT  15.90 2.40 16.50 3.00 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        LAYER metal1 ;
        RECT  8.70 17.70 9.90 24.90 ;
        RECT  8.70 2.10 9.90 7.80 ;
        RECT  0.60 8.40 6.60 9.60 ;
        RECT  12.00 14.70 13.20 15.90 ;
        RECT  0.60 15.00 13.20 15.90 ;
        RECT  0.60 2.10 1.80 24.90 ;
        RECT  2.70 10.50 13.20 11.40 ;
        RECT  2.70 10.50 3.90 11.70 ;
        RECT  12.00 10.50 13.20 11.70 ;
        RECT  13.50 8.10 14.70 9.30 ;
        LAYER via ;
        RECT  9.00 24.00 9.60 24.60 ;
        RECT  9.00 22.50 9.60 23.10 ;
        RECT  9.00 21.00 9.60 21.60 ;
        RECT  9.00 19.50 9.60 20.10 ;
        RECT  9.00 18.00 9.60 18.60 ;
        RECT  9.00 6.90 9.60 7.50 ;
        RECT  9.00 5.40 9.60 6.00 ;
        RECT  9.00 3.90 9.60 4.50 ;
        RECT  9.00 2.40 9.60 3.00 ;
        RECT  13.80 8.40 14.40 9.00 ;
        LAYER metal2 ;
        RECT  8.70 8.10 14.70 9.30 ;
        RECT  8.70 2.10 9.90 24.90 ;
    END
END MUX2X2

MACRO MUX2NX1
    CLASS CORE ;
    FOREIGN MUX2NX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 13.20 6.30 13.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 14.10 ;
        LAYER metal1 ;
        RECT  5.40 12.90 6.60 14.10 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  12.90 12.90 13.50 13.50 ;
        LAYER metal2 ;
        RECT  12.60 12.60 13.80 17.10 ;
        LAYER metal1 ;
        RECT  9.60 12.60 13.80 13.80 ;
        END
    END B
    PIN S
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.20 3.90 13.80 ;
        LAYER metal2 ;
        RECT  3.00 12.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 12.90 4.20 14.10 ;
        END
    END S
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  9.00 2.40 9.60 3.00 ;
        RECT  9.00 3.90 9.60 4.50 ;
        RECT  9.00 5.40 9.60 6.00 ;
        RECT  9.00 6.90 9.60 7.50 ;
        RECT  9.00 18.00 9.60 18.60 ;
        RECT  9.00 19.50 9.60 20.10 ;
        RECT  9.00 21.00 9.60 21.60 ;
        RECT  9.00 22.50 9.60 23.10 ;
        RECT  9.00 24.00 9.60 24.60 ;
        LAYER metal2 ;
        RECT  8.70 2.10 9.90 24.90 ;
        RECT  7.80 6.90 9.90 8.10 ;
        LAYER metal1 ;
        RECT  8.70 2.10 9.90 7.80 ;
        RECT  8.70 17.70 9.90 24.90 ;
        END
    END Y
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 15.60 1.20 ;
        RECT  12.60 -1.20 13.80 7.50 ;
        RECT  3.00 -1.20 5.70 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 15.60 28.20 ;
        RECT  12.60 18.00 13.80 28.20 ;
        RECT  3.00 18.00 5.70 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.00 10.80 3.60 11.40 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 13.20 3.90 13.80 ;
        RECT  3.30 6.60 3.90 7.20 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 24.30 5.40 24.90 ;
        RECT  4.80 22.80 5.40 23.40 ;
        RECT  4.80 21.30 5.40 21.90 ;
        RECT  4.80 19.80 5.40 20.40 ;
        RECT  4.80 18.30 5.40 18.90 ;
        RECT  4.80 6.60 5.40 7.20 ;
        RECT  4.80 5.10 5.40 5.70 ;
        RECT  4.80 3.60 5.40 4.20 ;
        RECT  4.80 2.10 5.40 2.70 ;
        RECT  5.40 8.70 6.00 9.30 ;
        RECT  5.70 13.20 6.30 13.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  9.00 24.00 9.60 24.60 ;
        RECT  9.00 22.50 9.60 23.10 ;
        RECT  9.00 21.00 9.60 21.60 ;
        RECT  9.00 19.50 9.60 20.10 ;
        RECT  9.00 18.00 9.60 18.60 ;
        RECT  9.00 6.90 9.60 7.50 ;
        RECT  9.00 5.40 9.60 6.00 ;
        RECT  9.00 3.90 9.60 4.50 ;
        RECT  9.00 2.40 9.60 3.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  9.90 12.90 10.50 13.50 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.30 15.00 12.90 15.60 ;
        RECT  12.30 10.80 12.90 11.40 ;
        RECT  12.90 24.30 13.50 24.90 ;
        RECT  12.90 22.80 13.50 23.40 ;
        RECT  12.90 21.30 13.50 21.90 ;
        RECT  12.90 19.80 13.50 20.40 ;
        RECT  12.90 18.30 13.50 18.90 ;
        RECT  12.90 6.60 13.50 7.20 ;
        RECT  12.90 5.10 13.50 5.70 ;
        RECT  12.90 3.60 13.50 4.20 ;
        RECT  12.90 2.10 13.50 2.70 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        LAYER metal1 ;
        RECT  0.60 8.40 6.60 9.60 ;
        RECT  12.00 14.70 13.20 15.90 ;
        RECT  0.60 15.00 13.20 15.90 ;
        RECT  0.60 2.10 1.80 24.90 ;
        RECT  2.70 10.50 13.20 11.40 ;
        RECT  2.70 10.50 3.90 11.70 ;
        RECT  12.00 10.50 13.20 11.70 ;
    END
END MUX2NX1

MACRO LCX1
    CLASS CORE ;
    FOREIGN LCX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 10.20 3.90 10.80 ;
        LAYER metal2 ;
        RECT  3.00 9.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 9.90 5.40 11.10 ;
        END
    END D
    PIN CLR
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  22.50 10.20 23.10 10.80 ;
        LAYER metal2 ;
        RECT  22.20 9.90 23.40 11.10 ;
        LAYER metal1 ;
        RECT  21.00 9.90 23.40 11.10 ;
        END
    END CLR
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  15.30 2.40 15.90 3.00 ;
        RECT  15.30 3.90 15.90 4.50 ;
        RECT  15.30 19.50 15.90 20.10 ;
        RECT  15.30 21.00 15.90 21.60 ;
        RECT  15.30 22.50 15.90 23.10 ;
        RECT  15.30 24.00 15.90 24.60 ;
        LAYER metal2 ;
        RECT  15.00 2.10 16.20 24.90 ;
        LAYER metal1 ;
        RECT  15.00 2.10 16.20 4.80 ;
        RECT  15.00 19.20 16.20 24.90 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  5.70 7.20 6.30 7.80 ;
        LAYER metal2 ;
        RECT  5.40 6.90 6.60 8.10 ;
        LAYER metal1 ;
        RECT  6.75 10.80 8.10 12.00 ;
        RECT  6.75 8.10 7.80 12.00 ;
        RECT  1.50 8.10 7.80 9.00 ;
        RECT  5.40 6.90 6.60 9.00 ;
        RECT  1.50 7.80 2.70 9.00 ;
        END
    END G
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 25.20 1.20 ;
        RECT  17.40 -1.20 18.60 7.50 ;
        RECT  12.60 -1.20 13.80 4.50 ;
        RECT  3.00 -1.20 4.20 6.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 25.20 28.20 ;
        RECT  22.20 19.50 23.40 28.20 ;
        RECT  17.40 19.50 18.60 28.20 ;
        RECT  12.60 18.00 13.80 28.20 ;
        RECT  3.00 18.00 4.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  1.80 8.10 2.40 8.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 10.20 5.10 10.80 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 15.00 7.80 15.60 ;
        RECT  7.20 11.10 7.80 11.70 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  9.00 8.40 9.60 9.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.40 12.90 12.00 13.50 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.90 24.30 13.50 24.90 ;
        RECT  12.90 22.80 13.50 23.40 ;
        RECT  12.90 21.30 13.50 21.90 ;
        RECT  12.90 19.80 13.50 20.40 ;
        RECT  12.90 18.30 13.50 18.90 ;
        RECT  12.90 3.60 13.50 4.20 ;
        RECT  12.90 2.10 13.50 2.70 ;
        RECT  13.80 12.90 14.40 13.50 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.30 24.00 15.90 24.60 ;
        RECT  15.30 22.50 15.90 23.10 ;
        RECT  15.30 21.00 15.90 21.60 ;
        RECT  15.30 19.50 15.90 20.10 ;
        RECT  15.30 3.90 15.90 4.50 ;
        RECT  15.30 2.40 15.90 3.00 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 24.30 18.30 24.90 ;
        RECT  17.70 22.80 18.30 23.40 ;
        RECT  17.70 21.30 18.30 21.90 ;
        RECT  17.70 19.80 18.30 20.40 ;
        RECT  17.70 8.70 18.30 9.30 ;
        RECT  17.70 6.60 18.30 7.20 ;
        RECT  17.70 5.10 18.30 5.70 ;
        RECT  17.70 3.60 18.30 4.20 ;
        RECT  17.70 2.10 18.30 2.70 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  20.10 24.00 20.70 24.60 ;
        RECT  20.10 22.50 20.70 23.10 ;
        RECT  20.10 21.00 20.70 21.60 ;
        RECT  20.10 19.50 20.70 20.10 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 10.20 21.90 10.80 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  21.60 6.90 22.20 7.50 ;
        RECT  21.60 5.40 22.20 6.00 ;
        RECT  21.60 3.90 22.20 4.50 ;
        RECT  21.60 2.40 22.20 3.00 ;
        RECT  22.50 24.30 23.10 24.90 ;
        RECT  22.50 22.80 23.10 23.40 ;
        RECT  22.50 21.30 23.10 21.90 ;
        RECT  22.50 19.80 23.10 20.40 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        LAYER metal1 ;
        RECT  0.60 19.20 1.80 24.90 ;
        RECT  0.60 2.10 1.80 4.80 ;
        RECT  7.80 17.70 9.00 24.90 ;
        RECT  7.80 2.10 9.00 4.80 ;
        RECT  8.70 8.10 9.90 9.30 ;
        RECT  9.00 8.10 9.90 15.90 ;
        RECT  0.60 14.70 9.90 15.90 ;
        RECT  7.80 5.70 16.35 6.90 ;
        RECT  15.15 5.70 16.35 9.45 ;
        RECT  15.15 8.40 18.60 9.45 ;
        RECT  17.40 8.40 18.60 9.60 ;
        RECT  19.80 19.20 21.00 24.90 ;
        RECT  11.10 12.60 21.00 13.80 ;
        RECT  21.30 2.10 22.50 7.80 ;
        RECT  19.80 5.10 22.50 7.80 ;
        LAYER via ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 15.00 1.50 15.60 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 6.00 8.70 6.60 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  20.10 24.00 20.70 24.60 ;
        RECT  20.10 22.50 20.70 23.10 ;
        RECT  20.10 21.00 20.70 21.60 ;
        RECT  20.10 19.50 20.70 20.10 ;
        RECT  20.10 12.90 20.70 13.50 ;
        RECT  20.10 6.90 20.70 7.50 ;
        RECT  20.10 5.40 20.70 6.00 ;
        LAYER metal2 ;
        RECT  0.60 2.10 1.80 24.90 ;
        RECT  7.80 2.10 9.00 24.90 ;
        RECT  19.80 5.10 21.00 24.90 ;
    END
END LCX1

MACRO LCNX1
    CLASS CORE ;
    FOREIGN LCNX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 24.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 10.20 3.90 10.80 ;
        LAYER metal2 ;
        RECT  3.00 9.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 9.90 5.70 11.10 ;
        END
    END D
    PIN CLR
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  22.50 10.20 23.10 10.80 ;
        LAYER metal2 ;
        RECT  22.20 9.90 23.40 11.10 ;
        LAYER metal1 ;
        RECT  21.00 9.90 23.40 11.10 ;
        END
    END CLR
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  15.30 2.40 15.90 3.00 ;
        RECT  15.30 3.90 15.90 4.50 ;
        RECT  15.30 19.50 15.90 20.10 ;
        RECT  15.30 21.00 15.90 21.60 ;
        RECT  15.30 22.50 15.90 23.10 ;
        RECT  15.30 24.00 15.90 24.60 ;
        LAYER metal2 ;
        RECT  15.00 2.10 16.20 24.90 ;
        LAYER metal1 ;
        RECT  15.00 2.10 16.20 4.80 ;
        RECT  15.00 19.20 16.20 24.90 ;
        END
    END Q
    PIN G
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  5.70 7.20 6.30 7.80 ;
        LAYER metal2 ;
        RECT  5.40 6.90 6.60 8.10 ;
        LAYER metal1 ;
        RECT  8.70 8.10 9.90 9.30 ;
        RECT  1.50 8.10 9.90 9.00 ;
        RECT  6.90 12.60 8.10 13.80 ;
        RECT  6.90 8.10 7.80 13.80 ;
        RECT  5.40 6.90 6.60 9.00 ;
        RECT  1.50 7.80 2.70 9.00 ;
        END
    END G
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 25.20 1.20 ;
        RECT  17.40 -1.20 18.60 7.50 ;
        RECT  12.60 -1.20 13.80 4.50 ;
        RECT  3.00 -1.20 4.20 6.00 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 25.20 28.20 ;
        RECT  22.20 19.50 23.40 28.20 ;
        RECT  17.40 19.50 18.60 28.20 ;
        RECT  12.60 18.00 13.80 28.20 ;
        RECT  3.00 18.00 4.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  1.80 8.10 2.40 8.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 10.20 5.40 10.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 12.90 7.80 13.50 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  9.00 15.00 9.60 15.60 ;
        RECT  9.00 8.40 9.60 9.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.40 12.90 12.00 13.50 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.90 24.30 13.50 24.90 ;
        RECT  12.90 22.80 13.50 23.40 ;
        RECT  12.90 21.30 13.50 21.90 ;
        RECT  12.90 19.80 13.50 20.40 ;
        RECT  12.90 18.30 13.50 18.90 ;
        RECT  12.90 3.60 13.50 4.20 ;
        RECT  12.90 2.10 13.50 2.70 ;
        RECT  13.80 12.90 14.40 13.50 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.30 24.00 15.90 24.60 ;
        RECT  15.30 22.50 15.90 23.10 ;
        RECT  15.30 21.00 15.90 21.60 ;
        RECT  15.30 19.50 15.90 20.10 ;
        RECT  15.30 3.90 15.90 4.50 ;
        RECT  15.30 2.40 15.90 3.00 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 24.30 18.30 24.90 ;
        RECT  17.70 22.80 18.30 23.40 ;
        RECT  17.70 21.30 18.30 21.90 ;
        RECT  17.70 19.80 18.30 20.40 ;
        RECT  17.70 8.70 18.30 9.30 ;
        RECT  17.70 6.60 18.30 7.20 ;
        RECT  17.70 5.10 18.30 5.70 ;
        RECT  17.70 3.60 18.30 4.20 ;
        RECT  17.70 2.10 18.30 2.70 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  20.10 24.00 20.70 24.60 ;
        RECT  20.10 22.50 20.70 23.10 ;
        RECT  20.10 21.00 20.70 21.60 ;
        RECT  20.10 19.50 20.70 20.10 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 10.20 21.90 10.80 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  21.60 6.90 22.20 7.50 ;
        RECT  21.60 5.40 22.20 6.00 ;
        RECT  21.60 3.90 22.20 4.50 ;
        RECT  21.60 2.40 22.20 3.00 ;
        RECT  22.50 24.30 23.10 24.90 ;
        RECT  22.50 22.80 23.10 23.40 ;
        RECT  22.50 21.30 23.10 21.90 ;
        RECT  22.50 19.80 23.10 20.40 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        LAYER metal1 ;
        RECT  0.60 19.20 1.80 24.90 ;
        RECT  0.60 2.10 1.80 4.80 ;
        RECT  7.80 17.70 9.00 24.90 ;
        RECT  7.80 2.10 9.00 4.80 ;
        RECT  0.60 14.70 1.80 15.90 ;
        RECT  8.70 14.70 9.90 15.90 ;
        RECT  0.60 15.00 9.90 15.90 ;
        RECT  7.80 5.70 16.35 6.90 ;
        RECT  15.15 5.70 16.35 9.45 ;
        RECT  15.15 8.40 18.60 9.45 ;
        RECT  17.40 8.40 18.60 9.60 ;
        RECT  19.80 19.20 21.00 24.90 ;
        RECT  11.10 12.60 21.00 13.80 ;
        RECT  21.30 2.10 22.50 7.80 ;
        RECT  19.80 5.10 22.50 7.80 ;
        LAYER via ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 15.00 1.50 15.60 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 6.00 8.70 6.60 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  20.10 24.00 20.70 24.60 ;
        RECT  20.10 22.50 20.70 23.10 ;
        RECT  20.10 21.00 20.70 21.60 ;
        RECT  20.10 19.50 20.70 20.10 ;
        RECT  20.10 12.90 20.70 13.50 ;
        RECT  20.10 6.90 20.70 7.50 ;
        RECT  20.10 5.40 20.70 6.00 ;
        LAYER metal2 ;
        RECT  0.60 2.10 1.80 24.90 ;
        RECT  7.80 2.10 9.00 24.90 ;
        RECT  19.80 5.10 21.00 24.90 ;
    END
END LCNX1

MACRO INVX8
    CLASS CORE ;
    FOREIGN INVX8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 13.50 8.70 14.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 24.00 8.70 24.60 ;
        LAYER metal2 ;
        RECT  7.80 2.10 9.00 24.90 ;
        LAYER metal1 ;
        RECT  7.80 2.10 9.00 24.90 ;
        RECT  3.00 11.70 9.00 12.60 ;
        RECT  3.00 8.40 9.00 9.30 ;
        RECT  3.00 2.10 4.20 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 13.20 28.20 ;
        RECT  10.20 13.50 11.40 28.20 ;
        RECT  5.40 13.50 6.60 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 13.20 1.20 ;
        RECT  10.20 -1.20 11.40 7.50 ;
        RECT  5.40 -1.20 6.60 7.50 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 18.30 6.30 18.90 ;
        RECT  5.70 16.80 6.30 17.40 ;
        RECT  5.70 15.30 6.30 15.90 ;
        RECT  5.70 13.80 6.30 14.40 ;
        RECT  5.70 6.60 6.30 7.20 ;
        RECT  5.70 5.10 6.30 5.70 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 13.50 8.70 14.10 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.50 24.30 11.10 24.90 ;
        RECT  10.50 22.80 11.10 23.40 ;
        RECT  10.50 21.30 11.10 21.90 ;
        RECT  10.50 19.80 11.10 20.40 ;
        RECT  10.50 18.30 11.10 18.90 ;
        RECT  10.50 16.80 11.10 17.40 ;
        RECT  10.50 15.30 11.10 15.90 ;
        RECT  10.50 13.80 11.10 14.40 ;
        RECT  10.50 6.60 11.10 7.20 ;
        RECT  10.50 5.10 11.10 5.70 ;
        RECT  10.50 3.60 11.10 4.20 ;
        RECT  10.50 2.10 11.10 2.70 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
    END
END INVX8

MACRO INVX4
    CLASS CORE ;
    FOREIGN INVX4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 24.90 ;
        LAYER metal1 ;
        RECT  3.00 2.10 4.20 7.80 ;
        RECT  3.00 13.20 4.20 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 8.40 28.20 ;
        RECT  5.40 13.50 6.60 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 8.40 1.20 ;
        RECT  5.40 -1.20 6.60 7.50 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 18.30 6.30 18.90 ;
        RECT  5.70 16.80 6.30 17.40 ;
        RECT  5.70 15.30 6.30 15.90 ;
        RECT  5.70 13.80 6.30 14.40 ;
        RECT  5.70 6.60 6.30 7.20 ;
        RECT  5.70 5.10 6.30 5.70 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
    END
END INVX4

MACRO INVX2
    CLASS CORE ;
    FOREIGN INVX2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        LAYER metal2 ;
        RECT  3.00 13.20 4.20 24.90 ;
        LAYER metal1 ;
        RECT  3.00 2.10 4.20 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 6.00 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 6.00 1.20 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
    END
END INVX2

MACRO INVX16
    CLASS CORE ;
    FOREIGN INVX16 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 21.60 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 13.50 8.70 14.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 24.00 8.70 24.60 ;
        LAYER metal2 ;
        RECT  7.80 2.10 9.00 24.90 ;
        LAYER metal1 ;
        RECT  17.40 2.10 18.60 24.90 ;
        RECT  3.00 11.70 18.60 12.60 ;
        RECT  3.00 8.40 18.60 9.30 ;
        RECT  12.60 2.10 13.80 24.90 ;
        RECT  7.80 2.10 9.00 24.90 ;
        RECT  3.00 2.10 4.20 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 22.80 28.20 ;
        RECT  19.80 13.50 21.00 28.20 ;
        RECT  15.00 13.50 16.20 28.20 ;
        RECT  10.20 13.50 11.40 28.20 ;
        RECT  5.40 13.50 6.60 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 22.80 1.20 ;
        RECT  19.80 -1.20 21.00 7.50 ;
        RECT  15.00 -1.20 16.20 7.50 ;
        RECT  10.20 -1.20 11.40 7.50 ;
        RECT  5.40 -1.20 6.60 7.50 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  8.10 13.50 8.70 14.10 ;
        RECT  10.50 24.30 11.10 24.90 ;
        RECT  10.50 22.80 11.10 23.40 ;
        RECT  10.50 21.30 11.10 21.90 ;
        RECT  10.50 19.80 11.10 20.40 ;
        RECT  10.50 18.30 11.10 18.90 ;
        RECT  10.50 16.80 11.10 17.40 ;
        RECT  10.50 15.30 11.10 15.90 ;
        RECT  10.50 13.80 11.10 14.40 ;
        RECT  10.50 6.60 11.10 7.20 ;
        RECT  10.50 5.10 11.10 5.70 ;
        RECT  10.50 3.60 11.10 4.20 ;
        RECT  10.50 2.10 11.10 2.70 ;
        RECT  12.90 13.50 13.50 14.10 ;
        RECT  17.70 13.50 18.30 14.10 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 6.60 6.30 7.20 ;
        RECT  5.70 5.10 6.30 5.70 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 18.30 6.30 18.90 ;
        RECT  5.70 16.80 6.30 17.40 ;
        RECT  5.70 15.30 6.30 15.90 ;
        RECT  5.70 13.80 6.30 14.40 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.90 6.90 13.50 7.50 ;
        RECT  12.90 5.40 13.50 6.00 ;
        RECT  12.90 3.90 13.50 4.50 ;
        RECT  12.90 2.40 13.50 3.00 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.30 6.60 15.90 7.20 ;
        RECT  15.30 5.10 15.90 5.70 ;
        RECT  15.30 3.60 15.90 4.20 ;
        RECT  15.30 2.10 15.90 2.70 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 6.90 18.30 7.50 ;
        RECT  17.70 5.40 18.30 6.00 ;
        RECT  17.70 3.90 18.30 4.50 ;
        RECT  17.70 2.40 18.30 3.00 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  20.10 6.60 20.70 7.20 ;
        RECT  20.10 5.10 20.70 5.70 ;
        RECT  20.10 3.60 20.70 4.20 ;
        RECT  20.10 2.10 20.70 2.70 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  12.90 24.00 13.50 24.60 ;
        RECT  12.90 22.50 13.50 23.10 ;
        RECT  12.90 21.00 13.50 21.60 ;
        RECT  12.90 19.50 13.50 20.10 ;
        RECT  12.90 18.00 13.50 18.60 ;
        RECT  12.90 16.50 13.50 17.10 ;
        RECT  12.90 15.00 13.50 15.60 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  15.30 24.30 15.90 24.90 ;
        RECT  15.30 22.80 15.90 23.40 ;
        RECT  15.30 21.30 15.90 21.90 ;
        RECT  15.30 19.80 15.90 20.40 ;
        RECT  15.30 18.30 15.90 18.90 ;
        RECT  15.30 16.80 15.90 17.40 ;
        RECT  15.30 15.30 15.90 15.90 ;
        RECT  15.30 13.80 15.90 14.40 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  17.70 24.00 18.30 24.60 ;
        RECT  17.70 22.50 18.30 23.10 ;
        RECT  17.70 21.00 18.30 21.60 ;
        RECT  17.70 19.50 18.30 20.10 ;
        RECT  17.70 18.00 18.30 18.60 ;
        RECT  17.70 16.50 18.30 17.10 ;
        RECT  17.70 15.00 18.30 15.60 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  20.10 24.30 20.70 24.90 ;
        RECT  20.10 22.80 20.70 23.40 ;
        RECT  20.10 21.30 20.70 21.90 ;
        RECT  20.10 19.80 20.70 20.40 ;
        RECT  20.10 18.30 20.70 18.90 ;
        RECT  20.10 16.80 20.70 17.40 ;
        RECT  20.10 15.30 20.70 15.90 ;
        RECT  20.10 13.80 20.70 14.40 ;
        RECT  21.30 26.70 21.90 27.30 ;
    END
END INVX16

MACRO INVX1
    CLASS CORE ;
    FOREIGN INVX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 4.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 16.20 3.90 16.80 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 24.90 ;
        LAYER metal1 ;
        RECT  3.00 2.10 4.20 4.80 ;
        RECT  3.00 15.90 4.20 17.10 ;
        RECT  3.00 19.20 4.20 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 6.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 6.00 1.20 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
    END
END INVX1

MACRO FILL8
    CLASS CORE ;
    FOREIGN FILL8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 36.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 37.20 1.20 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 37.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        RECT  26.10 26.70 26.70 27.30 ;
        RECT  26.10 -0.30 26.70 0.30 ;
        RECT  28.50 26.70 29.10 27.30 ;
        RECT  28.50 -0.30 29.10 0.30 ;
        RECT  30.90 26.70 31.50 27.30 ;
        RECT  30.90 -0.30 31.50 0.30 ;
        RECT  33.30 26.70 33.90 27.30 ;
        RECT  33.30 -0.30 33.90 0.30 ;
        RECT  35.70 26.70 36.30 27.30 ;
        RECT  35.70 -0.30 36.30 0.30 ;
    END
END FILL8

MACRO FILL4
    CLASS CORE ;
    FOREIGN FILL4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 18.00 1.20 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 18.00 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
    END
END FILL4

MACRO FILL2
    CLASS CORE ;
    FOREIGN FILL2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 8.40 1.20 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 8.40 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
    END
END FILL2

MACRO FILL
    CLASS CORE ;
    FOREIGN FILL 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 2.40 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 3.60 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 3.60 1.20 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
    END
END FILL

MACRO ENINVX2
    CLASS CORE ;
    FOREIGN ENINVX2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 14.40 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 2.55 1.50 3.15 ;
        LAYER metal2 ;
        RECT  0.60 2.25 1.80 5.10 ;
        LAYER metal1 ;
        RECT  0.60 2.25 3.00 3.45 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 24.00 8.70 24.60 ;
        LAYER metal2 ;
        RECT  7.80 3.60 9.00 25.20 ;
        LAYER metal1 ;
        RECT  7.80 3.60 9.00 7.80 ;
        RECT  7.80 14.70 9.00 24.90 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 10.20 6.30 10.80 ;
        LAYER metal2 ;
        RECT  5.40 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  5.40 9.90 11.85 11.10 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 15.60 1.20 ;
        RECT  11.70 -1.20 12.90 7.35 ;
        RECT  3.90 -1.20 5.10 7.35 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 15.60 28.20 ;
        RECT  11.70 14.70 12.90 28.20 ;
        RECT  3.90 14.70 5.10 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  1.80 24.00 2.40 24.60 ;
        RECT  1.80 22.50 2.40 23.10 ;
        RECT  1.80 21.00 2.40 21.60 ;
        RECT  1.80 19.50 2.40 20.10 ;
        RECT  1.80 6.45 2.40 7.05 ;
        RECT  1.80 4.95 2.40 5.55 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 2.55 2.70 3.15 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  4.20 24.00 4.80 24.60 ;
        RECT  4.20 22.50 4.80 23.10 ;
        RECT  4.20 21.00 4.80 21.60 ;
        RECT  4.20 19.50 4.80 20.10 ;
        RECT  4.20 18.00 4.80 18.60 ;
        RECT  4.20 16.50 4.80 17.10 ;
        RECT  4.20 15.00 4.80 15.60 ;
        RECT  4.20 6.45 4.80 7.05 ;
        RECT  4.20 4.95 4.80 5.55 ;
        RECT  4.20 3.45 4.80 4.05 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 10.20 6.30 10.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 12.30 8.70 12.90 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.95 10.20 11.55 10.80 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.00 24.00 12.60 24.60 ;
        RECT  12.00 22.50 12.60 23.10 ;
        RECT  12.00 21.00 12.60 21.60 ;
        RECT  12.00 19.50 12.60 20.10 ;
        RECT  12.00 18.00 12.60 18.60 ;
        RECT  12.00 16.50 12.60 17.10 ;
        RECT  12.00 15.00 12.60 15.60 ;
        RECT  12.00 6.45 12.60 7.05 ;
        RECT  12.00 4.95 12.60 5.55 ;
        RECT  12.00 3.45 12.60 4.05 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        LAYER metal1 ;
        RECT  1.50 12.00 9.00 13.20 ;
        RECT  1.50 4.65 2.70 24.90 ;
    END
END ENINVX2

MACRO ENINVX1
    CLASS CORE ;
    FOREIGN ENINVX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN EN
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 2.55 1.50 3.15 ;
        LAYER metal2 ;
        RECT  0.60 2.25 1.80 5.10 ;
        LAYER metal1 ;
        RECT  0.60 2.25 3.00 3.45 ;
        END
    END EN
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 24.00 8.70 24.60 ;
        LAYER metal2 ;
        RECT  7.80 3.60 9.00 25.20 ;
        LAYER metal1 ;
        RECT  7.80 3.60 9.00 7.80 ;
        RECT  7.80 14.70 9.00 24.90 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  4.80 10.20 5.40 10.80 ;
        LAYER metal2 ;
        RECT  4.50 9.90 6.60 11.10 ;
        LAYER metal1 ;
        RECT  4.50 9.90 5.70 11.10 ;
        END
    END A
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 10.80 1.20 ;
        RECT  3.90 -1.20 5.10 7.35 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 10.80 28.20 ;
        RECT  3.90 14.70 5.10 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  1.80 24.00 2.40 24.60 ;
        RECT  1.80 22.50 2.40 23.10 ;
        RECT  1.80 21.00 2.40 21.60 ;
        RECT  1.80 19.50 2.40 20.10 ;
        RECT  1.80 6.45 2.40 7.05 ;
        RECT  1.80 4.95 2.40 5.55 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 2.55 2.70 3.15 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  4.20 24.00 4.80 24.60 ;
        RECT  4.20 22.50 4.80 23.10 ;
        RECT  4.20 21.00 4.80 21.60 ;
        RECT  4.20 19.50 4.80 20.10 ;
        RECT  4.20 18.00 4.80 18.60 ;
        RECT  4.20 16.50 4.80 17.10 ;
        RECT  4.20 15.00 4.80 15.60 ;
        RECT  4.20 6.45 4.80 7.05 ;
        RECT  4.20 4.95 4.80 5.55 ;
        RECT  4.20 3.45 4.80 4.05 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  4.80 10.20 5.40 10.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 12.30 8.70 12.90 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        LAYER metal1 ;
        RECT  1.50 12.00 9.00 13.20 ;
        RECT  1.50 4.65 2.70 24.90 ;
    END
END ENINVX1

MACRO DCX1
    CLASS CORE ;
    FOREIGN DCX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 14.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 9.90 11.10 ;
        END
    END D
    PIN CLR
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  15.30 10.20 15.90 10.80 ;
        LAYER metal2 ;
        RECT  15.00 9.90 16.20 11.10 ;
        LAYER metal1 ;
        RECT  15.00 9.90 18.60 11.10 ;
        END
    END CLR
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  36.90 3.90 37.50 4.50 ;
        LAYER metal2 ;
        RECT  39.00 3.90 40.20 24.90 ;
        RECT  36.60 3.90 40.20 5.10 ;
        RECT  36.60 2.10 37.80 5.10 ;
        LAYER metal1 ;
        RECT  39.00 13.20 40.20 24.90 ;
        RECT  33.30 14.70 40.20 15.60 ;
        RECT  33.30 14.70 34.50 15.90 ;
        RECT  36.60 2.10 37.80 4.80 ;
        END
    END Q
    PIN CLK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 17.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 42.00 28.20 ;
        RECT  34.80 18.00 36.00 28.20 ;
        RECT  24.90 18.00 26.10 28.20 ;
        RECT  16.20 18.00 17.40 28.20 ;
        RECT  7.80 18.00 9.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 42.00 1.20 ;
        RECT  39.00 -1.20 40.20 4.50 ;
        RECT  34.20 -1.20 35.40 4.50 ;
        RECT  25.80 -1.20 27.00 6.00 ;
        RECT  21.00 -1.20 22.20 4.50 ;
        RECT  16.20 -1.20 17.40 4.50 ;
        RECT  7.80 -1.20 9.00 6.00 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  8.10 5.10 8.70 5.70 ;
        RECT  8.10 3.60 8.70 4.20 ;
        RECT  8.10 2.10 8.70 2.70 ;
        RECT  9.00 10.20 9.60 10.80 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.40 12.90 12.00 13.50 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  13.20 8.40 13.80 9.00 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.60 12.90 16.20 13.50 ;
        RECT  16.50 3.60 17.10 4.20 ;
        RECT  16.50 2.10 17.10 2.70 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 10.20 18.30 10.80 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  8.10 24.30 8.70 24.90 ;
        RECT  8.10 22.80 8.70 23.40 ;
        RECT  8.10 21.30 8.70 21.90 ;
        RECT  8.10 19.80 8.70 20.40 ;
        RECT  8.10 18.30 8.70 18.90 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  13.20 15.00 13.80 15.60 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 24.30 17.10 24.90 ;
        RECT  16.50 22.80 17.10 23.40 ;
        RECT  16.50 21.30 17.10 21.90 ;
        RECT  16.50 19.80 17.10 20.40 ;
        RECT  16.50 18.30 17.10 18.90 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  7.20 15.00 7.80 15.60 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  21.30 3.60 21.90 4.20 ;
        RECT  21.30 2.10 21.90 2.70 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  22.20 6.00 22.80 6.60 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        RECT  24.90 10.50 25.50 11.10 ;
        RECT  26.10 5.10 26.70 5.70 ;
        RECT  26.10 3.60 26.70 4.20 ;
        RECT  26.10 2.10 26.70 2.70 ;
        RECT  26.10 -0.30 26.70 0.30 ;
        RECT  27.00 12.60 27.60 13.20 ;
        RECT  28.50 -0.30 29.10 0.30 ;
        RECT  29.40 8.40 30.00 9.00 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  30.90 -0.30 31.50 0.30 ;
        RECT  31.20 12.90 31.80 13.50 ;
        RECT  33.30 -0.30 33.90 0.30 ;
        RECT  34.50 3.60 35.10 4.20 ;
        RECT  34.50 2.10 35.10 2.70 ;
        RECT  35.70 -0.30 36.30 0.30 ;
        RECT  36.00 10.50 36.60 11.10 ;
        RECT  36.90 3.90 37.50 4.50 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  37.80 6.00 38.40 6.60 ;
        RECT  38.10 -0.30 38.70 0.30 ;
        RECT  39.30 3.60 39.90 4.20 ;
        RECT  39.30 2.10 39.90 2.70 ;
        RECT  40.50 -0.30 41.10 0.30 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  25.20 24.30 25.80 24.90 ;
        RECT  25.20 22.80 25.80 23.40 ;
        RECT  25.20 21.30 25.80 21.90 ;
        RECT  25.20 19.80 25.80 20.40 ;
        RECT  25.20 18.30 25.80 18.90 ;
        RECT  26.10 26.70 26.70 27.30 ;
        RECT  28.50 26.70 29.10 27.30 ;
        RECT  29.40 15.00 30.00 15.60 ;
        RECT  30.30 24.00 30.90 24.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.90 26.70 31.50 27.30 ;
        RECT  33.30 26.70 33.90 27.30 ;
        RECT  33.60 15.00 34.20 15.60 ;
        RECT  35.10 24.30 35.70 24.90 ;
        RECT  35.10 22.80 35.70 23.40 ;
        RECT  35.10 21.30 35.70 21.90 ;
        RECT  35.10 19.80 35.70 20.40 ;
        RECT  35.10 18.30 35.70 18.90 ;
        RECT  35.70 26.70 36.30 27.30 ;
        RECT  38.10 26.70 38.70 27.30 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  40.50 26.70 41.10 27.30 ;
        LAYER metal1 ;
        RECT  3.00 19.20 4.20 24.90 ;
        RECT  3.00 2.10 4.20 4.80 ;
        RECT  5.40 19.20 6.60 24.90 ;
        RECT  5.40 2.10 6.60 4.80 ;
        RECT  12.00 17.70 13.20 24.90 ;
        RECT  12.00 2.10 13.20 4.80 ;
        RECT  18.60 19.20 19.80 24.90 ;
        RECT  18.60 2.10 19.80 4.80 ;
        RECT  21.00 17.70 22.20 24.90 ;
        RECT  12.00 5.70 23.10 6.60 ;
        RECT  12.00 5.70 13.20 6.90 ;
        RECT  21.90 5.70 23.10 6.90 ;
        RECT  23.40 2.10 24.60 4.80 ;
        RECT  26.70 12.30 27.90 13.50 ;
        RECT  15.30 12.60 27.90 13.50 ;
        RECT  15.30 12.60 16.50 13.80 ;
        RECT  21.00 12.60 22.20 13.80 ;
        RECT  23.40 12.60 24.60 13.80 ;
        RECT  3.00 14.70 8.10 15.90 ;
        RECT  12.90 14.70 14.10 15.90 ;
        RECT  29.10 14.70 30.30 15.90 ;
        RECT  3.00 15.00 30.30 15.90 ;
        RECT  30.00 17.70 31.20 24.90 ;
        RECT  30.90 12.60 33.30 13.80 ;
        RECT  5.40 8.10 33.45 9.00 ;
        RECT  5.40 8.10 6.60 9.30 ;
        RECT  12.90 8.10 14.10 9.30 ;
        RECT  29.10 8.10 30.30 9.30 ;
        RECT  32.25 8.10 33.45 9.30 ;
        RECT  11.10 8.10 12.00 13.80 ;
        RECT  11.10 12.60 12.30 13.80 ;
        RECT  19.50 10.20 20.70 11.40 ;
        RECT  24.60 10.20 25.80 11.40 ;
        RECT  35.70 10.20 36.90 11.40 ;
        RECT  19.50 10.50 36.90 11.40 ;
        RECT  30.00 2.10 31.20 6.90 ;
        RECT  37.50 5.70 38.70 6.90 ;
        RECT  30.00 6.00 38.70 6.90 ;
        LAYER via ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 8.40 6.30 9.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  12.30 6.00 12.90 6.60 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  19.80 10.50 20.40 11.10 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  21.30 12.90 21.90 13.50 ;
        RECT  23.70 12.90 24.30 13.50 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  30.30 24.00 30.90 24.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  32.40 12.90 33.00 13.50 ;
        RECT  32.55 8.40 33.15 9.00 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 24.90 ;
        RECT  5.40 2.10 6.60 24.90 ;
        RECT  12.00 2.10 13.20 24.90 ;
        RECT  18.60 10.20 20.70 11.40 ;
        RECT  18.60 2.10 19.80 24.90 ;
        RECT  23.40 2.10 24.60 13.80 ;
        RECT  21.00 12.60 24.60 13.80 ;
        RECT  21.00 12.60 22.20 24.90 ;
        RECT  30.00 2.10 31.20 24.90 ;
        RECT  32.25 8.10 33.45 13.80 ;
        RECT  32.10 12.60 33.45 13.80 ;
    END
END DCX1

MACRO DCNX1
    CLASS CORE ;
    FOREIGN DCNX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 14.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 9.90 11.10 ;
        END
    END D
    PIN CLR
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  15.30 10.20 15.90 10.80 ;
        LAYER metal2 ;
        RECT  15.00 9.90 16.20 11.10 ;
        LAYER metal1 ;
        RECT  15.00 9.90 18.60 11.10 ;
        END
    END CLR
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  36.90 3.90 37.50 4.50 ;
        LAYER metal2 ;
        RECT  39.00 3.90 40.20 24.90 ;
        RECT  36.60 3.90 40.20 5.10 ;
        RECT  36.60 2.10 37.80 5.10 ;
        LAYER metal1 ;
        RECT  39.00 13.20 40.20 24.90 ;
        RECT  33.30 14.70 40.20 15.60 ;
        RECT  33.30 14.70 34.50 15.90 ;
        RECT  36.60 2.10 37.80 4.80 ;
        END
    END Q
    PIN CLK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 17.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END CLK
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 42.00 28.20 ;
        RECT  34.80 18.00 36.00 28.20 ;
        RECT  24.90 18.00 26.10 28.20 ;
        RECT  16.20 18.00 17.40 28.20 ;
        RECT  7.80 18.00 9.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 42.00 1.20 ;
        RECT  39.00 -1.20 40.20 4.50 ;
        RECT  34.20 -1.20 35.40 4.50 ;
        RECT  25.80 -1.20 27.00 6.00 ;
        RECT  21.00 -1.20 22.20 4.50 ;
        RECT  16.20 -1.20 17.40 4.50 ;
        RECT  7.80 -1.20 9.00 6.00 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  8.10 5.10 8.70 5.70 ;
        RECT  8.10 3.60 8.70 4.20 ;
        RECT  8.10 2.10 8.70 2.70 ;
        RECT  9.00 10.20 9.60 10.80 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.40 12.90 12.00 13.50 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  13.20 8.40 13.80 9.00 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.60 12.90 16.20 13.50 ;
        RECT  16.50 3.60 17.10 4.20 ;
        RECT  16.50 2.10 17.10 2.70 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 10.20 18.30 10.80 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  6.60 8.10 7.20 8.70 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  8.10 24.30 8.70 24.90 ;
        RECT  8.10 22.80 8.70 23.40 ;
        RECT  8.10 21.30 8.70 21.90 ;
        RECT  8.10 19.80 8.70 20.40 ;
        RECT  8.10 18.30 8.70 18.90 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  13.20 15.00 13.80 15.60 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 24.30 17.10 24.90 ;
        RECT  16.50 22.80 17.10 23.40 ;
        RECT  16.50 21.30 17.10 21.90 ;
        RECT  16.50 19.80 17.10 20.40 ;
        RECT  16.50 18.30 17.10 18.90 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  21.30 3.60 21.90 4.20 ;
        RECT  21.30 2.10 21.90 2.70 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  22.20 6.00 22.80 6.60 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        RECT  24.90 10.50 25.50 11.10 ;
        RECT  26.10 5.10 26.70 5.70 ;
        RECT  26.10 3.60 26.70 4.20 ;
        RECT  26.10 2.10 26.70 2.70 ;
        RECT  26.10 -0.30 26.70 0.30 ;
        RECT  27.00 12.60 27.60 13.20 ;
        RECT  28.50 -0.30 29.10 0.30 ;
        RECT  29.40 8.40 30.00 9.00 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  30.90 -0.30 31.50 0.30 ;
        RECT  31.20 12.90 31.80 13.50 ;
        RECT  33.30 -0.30 33.90 0.30 ;
        RECT  34.50 3.60 35.10 4.20 ;
        RECT  34.50 2.10 35.10 2.70 ;
        RECT  35.70 -0.30 36.30 0.30 ;
        RECT  36.00 10.50 36.60 11.10 ;
        RECT  36.90 3.90 37.50 4.50 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  37.80 6.00 38.40 6.60 ;
        RECT  38.10 -0.30 38.70 0.30 ;
        RECT  39.30 3.60 39.90 4.20 ;
        RECT  39.30 2.10 39.90 2.70 ;
        RECT  40.50 -0.30 41.10 0.30 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  25.20 24.30 25.80 24.90 ;
        RECT  25.20 22.80 25.80 23.40 ;
        RECT  25.20 21.30 25.80 21.90 ;
        RECT  25.20 19.80 25.80 20.40 ;
        RECT  25.20 18.30 25.80 18.90 ;
        RECT  26.10 26.70 26.70 27.30 ;
        RECT  28.50 26.70 29.10 27.30 ;
        RECT  29.40 15.00 30.00 15.60 ;
        RECT  30.30 24.00 30.90 24.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.90 26.70 31.50 27.30 ;
        RECT  33.30 26.70 33.90 27.30 ;
        RECT  33.60 15.00 34.20 15.60 ;
        RECT  35.10 24.30 35.70 24.90 ;
        RECT  35.10 22.80 35.70 23.40 ;
        RECT  35.10 21.30 35.70 21.90 ;
        RECT  35.10 19.80 35.70 20.40 ;
        RECT  35.10 18.30 35.70 18.90 ;
        RECT  35.70 26.70 36.30 27.30 ;
        RECT  38.10 26.70 38.70 27.30 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  40.50 26.70 41.10 27.30 ;
        LAYER metal1 ;
        RECT  3.00 19.20 4.20 24.90 ;
        RECT  3.00 2.10 4.20 4.80 ;
        RECT  5.40 19.20 6.60 24.90 ;
        RECT  5.40 2.10 6.60 4.80 ;
        RECT  12.00 17.70 13.20 24.90 ;
        RECT  12.00 2.10 13.20 4.80 ;
        RECT  18.60 19.20 19.80 24.90 ;
        RECT  18.60 2.10 19.80 4.80 ;
        RECT  21.00 17.70 22.20 24.90 ;
        RECT  12.00 5.70 23.10 6.60 ;
        RECT  12.00 5.70 13.20 6.90 ;
        RECT  21.90 5.70 23.10 6.90 ;
        RECT  23.40 2.10 24.60 4.80 ;
        RECT  26.70 12.30 27.90 13.50 ;
        RECT  15.30 12.60 27.90 13.50 ;
        RECT  15.30 12.60 16.50 13.80 ;
        RECT  21.00 12.60 22.20 13.80 ;
        RECT  23.40 12.60 24.60 13.80 ;
        RECT  5.40 14.70 6.60 15.90 ;
        RECT  12.90 14.70 14.10 15.90 ;
        RECT  29.10 14.70 30.30 15.90 ;
        RECT  5.40 15.00 30.30 15.90 ;
        RECT  30.00 17.70 31.20 24.90 ;
        RECT  30.90 12.60 33.30 13.80 ;
        RECT  6.30 7.80 7.50 9.00 ;
        RECT  3.00 8.10 33.45 9.00 ;
        RECT  3.00 8.10 4.20 9.30 ;
        RECT  12.90 8.10 14.10 9.30 ;
        RECT  29.10 8.10 30.30 9.30 ;
        RECT  32.25 8.10 33.45 9.30 ;
        RECT  11.10 8.10 12.00 13.80 ;
        RECT  11.10 12.60 12.30 13.80 ;
        RECT  19.50 10.20 20.70 11.40 ;
        RECT  24.60 10.20 25.80 11.40 ;
        RECT  35.70 10.20 36.90 11.40 ;
        RECT  19.50 10.50 36.90 11.40 ;
        RECT  30.00 2.10 31.20 6.90 ;
        RECT  37.50 5.70 38.70 6.90 ;
        RECT  30.00 6.00 38.70 6.90 ;
        LAYER via ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 8.40 3.90 9.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  12.30 6.00 12.90 6.60 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  19.80 10.50 20.40 11.10 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  21.30 12.90 21.90 13.50 ;
        RECT  23.70 12.90 24.30 13.50 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  30.30 24.00 30.90 24.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  32.40 12.90 33.00 13.50 ;
        RECT  32.55 8.40 33.15 9.00 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 24.90 ;
        RECT  5.40 2.10 6.60 24.90 ;
        RECT  12.00 2.10 13.20 24.90 ;
        RECT  18.60 10.20 20.70 11.40 ;
        RECT  18.60 2.10 19.80 24.90 ;
        RECT  23.40 2.10 24.60 13.80 ;
        RECT  21.00 12.60 24.60 13.80 ;
        RECT  21.00 12.60 22.20 24.90 ;
        RECT  30.00 2.10 31.20 24.90 ;
        RECT  32.25 8.10 33.45 13.80 ;
        RECT  32.10 12.60 33.45 13.80 ;
    END
END DCNX1

MACRO DCBX1
    CLASS CORE ;
    FOREIGN DCBX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 14.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 9.90 11.10 ;
        END
    END D
    PIN CLR
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  15.30 10.20 15.90 10.80 ;
        LAYER metal2 ;
        RECT  15.00 9.90 16.20 11.10 ;
        LAYER metal1 ;
        RECT  15.00 9.90 18.60 11.10 ;
        END
    END CLR
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  36.90 3.90 37.50 4.50 ;
        LAYER metal2 ;
        RECT  39.00 3.90 40.20 24.90 ;
        RECT  36.60 3.90 40.20 5.10 ;
        RECT  36.60 2.10 37.80 5.10 ;
        LAYER metal1 ;
        RECT  39.00 13.20 40.20 24.90 ;
        RECT  33.30 14.70 40.20 15.60 ;
        RECT  33.30 14.70 34.50 15.90 ;
        RECT  36.60 2.10 37.80 4.80 ;
        END
    END Q
    PIN CLK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 17.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END CLK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 24.00 30.90 24.60 ;
        LAYER metal2 ;
        RECT  30.00 2.10 31.20 24.90 ;
        RECT  29.40 6.90 31.20 8.10 ;
        LAYER metal1 ;
        RECT  30.00 6.00 38.70 6.90 ;
        RECT  37.50 5.70 38.70 6.90 ;
        RECT  30.00 2.10 31.20 6.90 ;
        RECT  30.00 17.70 31.20 24.90 ;
        END
    END QB
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 42.00 28.20 ;
        RECT  34.80 18.00 36.00 28.20 ;
        RECT  24.90 18.00 26.10 28.20 ;
        RECT  16.20 18.00 17.40 28.20 ;
        RECT  7.80 18.00 9.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 42.00 1.20 ;
        RECT  39.00 -1.20 40.20 4.50 ;
        RECT  34.20 -1.20 35.40 4.50 ;
        RECT  25.80 -1.20 27.00 6.00 ;
        RECT  21.00 -1.20 22.20 4.50 ;
        RECT  16.20 -1.20 17.40 4.50 ;
        RECT  7.80 -1.20 9.00 6.00 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  8.10 5.10 8.70 5.70 ;
        RECT  8.10 3.60 8.70 4.20 ;
        RECT  8.10 2.10 8.70 2.70 ;
        RECT  9.00 10.20 9.60 10.80 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.40 12.90 12.00 13.50 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  13.20 8.40 13.80 9.00 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.60 12.90 16.20 13.50 ;
        RECT  16.50 3.60 17.10 4.20 ;
        RECT  16.50 2.10 17.10 2.70 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 10.20 18.30 10.80 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  8.10 24.30 8.70 24.90 ;
        RECT  8.10 22.80 8.70 23.40 ;
        RECT  8.10 21.30 8.70 21.90 ;
        RECT  8.10 19.80 8.70 20.40 ;
        RECT  8.10 18.30 8.70 18.90 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  13.20 15.00 13.80 15.60 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 24.30 17.10 24.90 ;
        RECT  16.50 22.80 17.10 23.40 ;
        RECT  16.50 21.30 17.10 21.90 ;
        RECT  16.50 19.80 17.10 20.40 ;
        RECT  16.50 18.30 17.10 18.90 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  7.20 15.00 7.80 15.60 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  21.30 3.60 21.90 4.20 ;
        RECT  21.30 2.10 21.90 2.70 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  22.20 6.00 22.80 6.60 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        RECT  24.90 10.50 25.50 11.10 ;
        RECT  26.10 5.10 26.70 5.70 ;
        RECT  26.10 3.60 26.70 4.20 ;
        RECT  26.10 2.10 26.70 2.70 ;
        RECT  26.10 -0.30 26.70 0.30 ;
        RECT  27.00 12.60 27.60 13.20 ;
        RECT  28.50 -0.30 29.10 0.30 ;
        RECT  29.40 8.40 30.00 9.00 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  30.90 -0.30 31.50 0.30 ;
        RECT  31.20 12.90 31.80 13.50 ;
        RECT  33.30 -0.30 33.90 0.30 ;
        RECT  34.50 3.60 35.10 4.20 ;
        RECT  34.50 2.10 35.10 2.70 ;
        RECT  35.70 -0.30 36.30 0.30 ;
        RECT  36.00 10.50 36.60 11.10 ;
        RECT  36.90 3.90 37.50 4.50 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  37.80 6.00 38.40 6.60 ;
        RECT  38.10 -0.30 38.70 0.30 ;
        RECT  39.30 3.60 39.90 4.20 ;
        RECT  39.30 2.10 39.90 2.70 ;
        RECT  40.50 -0.30 41.10 0.30 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  25.20 24.30 25.80 24.90 ;
        RECT  25.20 22.80 25.80 23.40 ;
        RECT  25.20 21.30 25.80 21.90 ;
        RECT  25.20 19.80 25.80 20.40 ;
        RECT  25.20 18.30 25.80 18.90 ;
        RECT  26.10 26.70 26.70 27.30 ;
        RECT  28.50 26.70 29.10 27.30 ;
        RECT  29.40 15.00 30.00 15.60 ;
        RECT  30.30 24.00 30.90 24.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.90 26.70 31.50 27.30 ;
        RECT  33.30 26.70 33.90 27.30 ;
        RECT  33.60 15.00 34.20 15.60 ;
        RECT  35.10 24.30 35.70 24.90 ;
        RECT  35.10 22.80 35.70 23.40 ;
        RECT  35.10 21.30 35.70 21.90 ;
        RECT  35.10 19.80 35.70 20.40 ;
        RECT  35.10 18.30 35.70 18.90 ;
        RECT  35.70 26.70 36.30 27.30 ;
        RECT  38.10 26.70 38.70 27.30 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  40.50 26.70 41.10 27.30 ;
        LAYER metal1 ;
        RECT  3.00 19.20 4.20 24.90 ;
        RECT  3.00 2.10 4.20 4.80 ;
        RECT  5.40 19.20 6.60 24.90 ;
        RECT  5.40 2.10 6.60 4.80 ;
        RECT  12.00 17.70 13.20 24.90 ;
        RECT  12.00 2.10 13.20 4.80 ;
        RECT  18.60 19.20 19.80 24.90 ;
        RECT  18.60 2.10 19.80 4.80 ;
        RECT  21.00 17.70 22.20 24.90 ;
        RECT  12.00 5.70 23.10 6.60 ;
        RECT  12.00 5.70 13.20 6.90 ;
        RECT  21.90 5.70 23.10 6.90 ;
        RECT  23.40 2.10 24.60 4.80 ;
        RECT  26.70 12.30 27.90 13.50 ;
        RECT  15.30 12.60 27.90 13.50 ;
        RECT  15.30 12.60 16.50 13.80 ;
        RECT  21.00 12.60 22.20 13.80 ;
        RECT  23.40 12.60 24.60 13.80 ;
        RECT  3.00 14.70 8.10 15.90 ;
        RECT  12.90 14.70 14.10 15.90 ;
        RECT  29.10 14.70 30.30 15.90 ;
        RECT  3.00 15.00 30.30 15.90 ;
        RECT  30.90 12.60 33.30 13.80 ;
        RECT  5.40 8.10 33.45 9.00 ;
        RECT  5.40 8.10 6.60 9.30 ;
        RECT  12.90 8.10 14.10 9.30 ;
        RECT  29.10 8.10 30.30 9.30 ;
        RECT  32.25 8.10 33.45 9.30 ;
        RECT  11.10 8.10 12.00 13.80 ;
        RECT  11.10 12.60 12.30 13.80 ;
        RECT  19.50 10.20 20.70 11.40 ;
        RECT  24.60 10.20 25.80 11.40 ;
        RECT  35.70 10.20 36.90 11.40 ;
        RECT  19.50 10.50 36.90 11.40 ;
        LAYER via ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 8.40 6.30 9.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  12.30 6.00 12.90 6.60 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  19.80 10.50 20.40 11.10 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  21.30 12.90 21.90 13.50 ;
        RECT  23.70 12.90 24.30 13.50 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  32.40 12.90 33.00 13.50 ;
        RECT  32.55 8.40 33.15 9.00 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 24.90 ;
        RECT  5.40 2.10 6.60 24.90 ;
        RECT  12.00 2.10 13.20 24.90 ;
        RECT  18.60 10.20 20.70 11.40 ;
        RECT  18.60 2.10 19.80 24.90 ;
        RECT  23.40 2.10 24.60 13.80 ;
        RECT  21.00 12.60 24.60 13.80 ;
        RECT  21.00 12.60 22.20 24.90 ;
        RECT  32.25 8.10 33.45 13.80 ;
        RECT  32.10 12.60 33.45 13.80 ;
    END
END DCBX1

MACRO DCBNX1
    CLASS CORE ;
    FOREIGN DCBNX1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 40.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 14.10 ;
        LAYER metal1 ;
        RECT  7.80 9.90 9.90 11.10 ;
        END
    END D
    PIN CLR
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  15.30 10.20 15.90 10.80 ;
        LAYER metal2 ;
        RECT  15.00 9.90 16.20 11.10 ;
        LAYER metal1 ;
        RECT  15.00 9.90 18.60 11.10 ;
        END
    END CLR
    PIN Q
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  36.90 3.90 37.50 4.50 ;
        LAYER metal2 ;
        RECT  39.00 3.90 40.20 24.90 ;
        RECT  36.60 3.90 40.20 5.10 ;
        RECT  36.60 2.10 37.80 5.10 ;
        LAYER metal1 ;
        RECT  39.00 13.20 40.20 24.90 ;
        RECT  33.30 14.70 40.20 15.60 ;
        RECT  33.30 14.70 34.50 15.90 ;
        RECT  36.60 2.10 37.80 4.80 ;
        END
    END Q
    PIN CLK
        DIRECTION INPUT ;
        USE CLOCK ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 17.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END CLK
    PIN QB
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 24.00 30.90 24.60 ;
        LAYER metal2 ;
        RECT  30.00 2.10 31.20 24.90 ;
        RECT  29.40 6.90 31.20 8.10 ;
        LAYER metal1 ;
        RECT  30.00 6.00 38.70 6.90 ;
        RECT  37.50 5.70 38.70 6.90 ;
        RECT  30.00 2.10 31.20 6.90 ;
        RECT  30.00 17.70 31.20 24.90 ;
        END
    END QB
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 42.00 28.20 ;
        RECT  34.80 18.00 36.00 28.20 ;
        RECT  24.90 18.00 26.10 28.20 ;
        RECT  16.20 18.00 17.40 28.20 ;
        RECT  7.80 18.00 9.00 28.20 ;
        RECT  0.60 19.50 1.80 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 42.00 1.20 ;
        RECT  39.00 -1.20 40.20 4.50 ;
        RECT  34.20 -1.20 35.40 4.50 ;
        RECT  25.80 -1.20 27.00 6.00 ;
        RECT  21.00 -1.20 22.20 4.50 ;
        RECT  16.20 -1.20 17.40 4.50 ;
        RECT  7.80 -1.20 9.00 6.00 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  8.10 5.10 8.70 5.70 ;
        RECT  8.10 3.60 8.70 4.20 ;
        RECT  8.10 2.10 8.70 2.70 ;
        RECT  9.00 10.20 9.60 10.80 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  11.40 12.90 12.00 13.50 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  13.20 8.40 13.80 9.00 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.60 12.90 16.20 13.50 ;
        RECT  16.50 3.60 17.10 4.20 ;
        RECT  16.50 2.10 17.10 2.70 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        RECT  17.70 10.20 18.30 10.80 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  18.90 -0.30 19.50 0.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  6.60 8.10 7.20 8.70 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  8.10 24.30 8.70 24.90 ;
        RECT  8.10 22.80 8.70 23.40 ;
        RECT  8.10 21.30 8.70 21.90 ;
        RECT  8.10 19.80 8.70 20.40 ;
        RECT  8.10 18.30 8.70 18.90 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  13.20 15.00 13.80 15.60 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 24.30 17.10 24.90 ;
        RECT  16.50 22.80 17.10 23.40 ;
        RECT  16.50 21.30 17.10 21.90 ;
        RECT  16.50 19.80 17.10 20.40 ;
        RECT  16.50 18.30 17.10 18.90 ;
        RECT  18.90 26.70 19.50 27.30 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  21.30 3.60 21.90 4.20 ;
        RECT  21.30 2.10 21.90 2.70 ;
        RECT  21.30 -0.30 21.90 0.30 ;
        RECT  22.20 6.00 22.80 6.60 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  23.70 -0.30 24.30 0.30 ;
        RECT  24.90 10.50 25.50 11.10 ;
        RECT  26.10 5.10 26.70 5.70 ;
        RECT  26.10 3.60 26.70 4.20 ;
        RECT  26.10 2.10 26.70 2.70 ;
        RECT  26.10 -0.30 26.70 0.30 ;
        RECT  27.00 12.60 27.60 13.20 ;
        RECT  28.50 -0.30 29.10 0.30 ;
        RECT  29.40 8.40 30.00 9.00 ;
        RECT  30.30 5.40 30.90 6.00 ;
        RECT  30.30 3.90 30.90 4.50 ;
        RECT  30.30 2.40 30.90 3.00 ;
        RECT  30.90 -0.30 31.50 0.30 ;
        RECT  31.20 12.90 31.80 13.50 ;
        RECT  33.30 -0.30 33.90 0.30 ;
        RECT  34.50 3.60 35.10 4.20 ;
        RECT  34.50 2.10 35.10 2.70 ;
        RECT  35.70 -0.30 36.30 0.30 ;
        RECT  36.00 10.50 36.60 11.10 ;
        RECT  36.90 3.90 37.50 4.50 ;
        RECT  36.90 2.40 37.50 3.00 ;
        RECT  37.80 6.00 38.40 6.60 ;
        RECT  38.10 -0.30 38.70 0.30 ;
        RECT  39.30 3.60 39.90 4.20 ;
        RECT  39.30 2.10 39.90 2.70 ;
        RECT  40.50 -0.30 41.10 0.30 ;
        RECT  21.30 26.70 21.90 27.30 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  23.70 26.70 24.30 27.30 ;
        RECT  25.20 24.30 25.80 24.90 ;
        RECT  25.20 22.80 25.80 23.40 ;
        RECT  25.20 21.30 25.80 21.90 ;
        RECT  25.20 19.80 25.80 20.40 ;
        RECT  25.20 18.30 25.80 18.90 ;
        RECT  26.10 26.70 26.70 27.30 ;
        RECT  28.50 26.70 29.10 27.30 ;
        RECT  29.40 15.00 30.00 15.60 ;
        RECT  30.30 24.00 30.90 24.60 ;
        RECT  30.30 22.50 30.90 23.10 ;
        RECT  30.30 21.00 30.90 21.60 ;
        RECT  30.30 19.50 30.90 20.10 ;
        RECT  30.30 18.00 30.90 18.60 ;
        RECT  30.90 26.70 31.50 27.30 ;
        RECT  33.30 26.70 33.90 27.30 ;
        RECT  33.60 15.00 34.20 15.60 ;
        RECT  35.10 24.30 35.70 24.90 ;
        RECT  35.10 22.80 35.70 23.40 ;
        RECT  35.10 21.30 35.70 21.90 ;
        RECT  35.10 19.80 35.70 20.40 ;
        RECT  35.10 18.30 35.70 18.90 ;
        RECT  35.70 26.70 36.30 27.30 ;
        RECT  38.10 26.70 38.70 27.30 ;
        RECT  39.30 24.00 39.90 24.60 ;
        RECT  39.30 22.50 39.90 23.10 ;
        RECT  39.30 21.00 39.90 21.60 ;
        RECT  39.30 19.50 39.90 20.10 ;
        RECT  39.30 18.00 39.90 18.60 ;
        RECT  39.30 16.50 39.90 17.10 ;
        RECT  39.30 15.00 39.90 15.60 ;
        RECT  40.50 26.70 41.10 27.30 ;
        LAYER metal1 ;
        RECT  3.00 19.20 4.20 24.90 ;
        RECT  3.00 2.10 4.20 4.80 ;
        RECT  5.40 19.20 6.60 24.90 ;
        RECT  5.40 2.10 6.60 4.80 ;
        RECT  12.00 17.70 13.20 24.90 ;
        RECT  12.00 2.10 13.20 4.80 ;
        RECT  18.60 19.20 19.80 24.90 ;
        RECT  18.60 2.10 19.80 4.80 ;
        RECT  21.00 17.70 22.20 24.90 ;
        RECT  12.00 5.70 23.10 6.60 ;
        RECT  12.00 5.70 13.20 6.90 ;
        RECT  21.90 5.70 23.10 6.90 ;
        RECT  23.40 2.10 24.60 4.80 ;
        RECT  26.70 12.30 27.90 13.50 ;
        RECT  15.30 12.60 27.90 13.50 ;
        RECT  15.30 12.60 16.50 13.80 ;
        RECT  21.00 12.60 22.20 13.80 ;
        RECT  23.40 12.60 24.60 13.80 ;
        RECT  5.40 14.70 6.60 15.90 ;
        RECT  12.90 14.70 14.10 15.90 ;
        RECT  29.10 14.70 30.30 15.90 ;
        RECT  5.40 15.00 30.30 15.90 ;
        RECT  30.90 12.60 33.30 13.80 ;
        RECT  6.30 7.80 7.50 9.00 ;
        RECT  3.00 8.10 33.45 9.00 ;
        RECT  3.00 8.10 4.20 9.30 ;
        RECT  12.90 8.10 14.10 9.30 ;
        RECT  29.10 8.10 30.30 9.30 ;
        RECT  32.25 8.10 33.45 9.30 ;
        RECT  11.10 8.10 12.00 13.80 ;
        RECT  11.10 12.60 12.30 13.80 ;
        RECT  19.50 10.20 20.70 11.40 ;
        RECT  24.60 10.20 25.80 11.40 ;
        RECT  35.70 10.20 36.90 11.40 ;
        RECT  19.50 10.50 36.90 11.40 ;
        LAYER via ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 8.40 3.90 9.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  12.30 24.00 12.90 24.60 ;
        RECT  12.30 22.50 12.90 23.10 ;
        RECT  12.30 21.00 12.90 21.60 ;
        RECT  12.30 19.50 12.90 20.10 ;
        RECT  12.30 18.00 12.90 18.60 ;
        RECT  12.30 6.00 12.90 6.60 ;
        RECT  12.30 3.90 12.90 4.50 ;
        RECT  12.30 2.40 12.90 3.00 ;
        RECT  18.90 24.00 19.50 24.60 ;
        RECT  18.90 22.50 19.50 23.10 ;
        RECT  18.90 21.00 19.50 21.60 ;
        RECT  18.90 19.50 19.50 20.10 ;
        RECT  18.90 3.90 19.50 4.50 ;
        RECT  18.90 2.40 19.50 3.00 ;
        RECT  19.80 10.50 20.40 11.10 ;
        RECT  21.30 24.00 21.90 24.60 ;
        RECT  21.30 22.50 21.90 23.10 ;
        RECT  21.30 21.00 21.90 21.60 ;
        RECT  21.30 19.50 21.90 20.10 ;
        RECT  21.30 18.00 21.90 18.60 ;
        RECT  21.30 12.90 21.90 13.50 ;
        RECT  23.70 12.90 24.30 13.50 ;
        RECT  23.70 3.90 24.30 4.50 ;
        RECT  23.70 2.40 24.30 3.00 ;
        RECT  32.40 12.90 33.00 13.50 ;
        RECT  32.55 8.40 33.15 9.00 ;
        LAYER metal2 ;
        RECT  3.00 2.10 4.20 24.90 ;
        RECT  5.40 2.10 6.60 24.90 ;
        RECT  12.00 2.10 13.20 24.90 ;
        RECT  18.60 10.20 20.70 11.40 ;
        RECT  18.60 2.10 19.80 24.90 ;
        RECT  23.40 2.10 24.60 13.80 ;
        RECT  21.00 12.60 24.60 13.80 ;
        RECT  21.00 12.60 22.20 24.90 ;
        RECT  32.25 8.10 33.45 13.80 ;
        RECT  32.10 12.60 33.45 13.80 ;
    END
END DCBNX1

MACRO BUFX8
    CLASS CORE ;
    FOREIGN BUFX8 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  12.90 2.40 13.50 3.00 ;
        RECT  12.90 3.90 13.50 4.50 ;
        RECT  12.90 5.40 13.50 6.00 ;
        RECT  12.90 6.90 13.50 7.50 ;
        RECT  12.90 13.50 13.50 14.10 ;
        RECT  12.90 15.00 13.50 15.60 ;
        RECT  12.90 16.50 13.50 17.10 ;
        RECT  12.90 18.00 13.50 18.60 ;
        RECT  12.90 19.50 13.50 20.10 ;
        RECT  12.90 21.00 13.50 21.60 ;
        RECT  12.90 22.50 13.50 23.10 ;
        RECT  12.90 24.00 13.50 24.60 ;
        LAYER metal2 ;
        RECT  12.60 2.10 13.80 24.90 ;
        LAYER metal1 ;
        RECT  12.60 2.10 13.80 24.90 ;
        RECT  7.80 11.70 13.80 12.60 ;
        RECT  7.80 8.40 13.80 9.30 ;
        RECT  7.80 2.10 9.00 24.90 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END A
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 18.00 1.20 ;
        RECT  15.00 -1.20 16.20 7.50 ;
        RECT  10.20 -1.20 11.40 7.50 ;
        RECT  5.40 -1.20 6.60 7.50 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 18.00 28.20 ;
        RECT  15.00 13.50 16.20 28.20 ;
        RECT  10.20 13.50 11.40 28.20 ;
        RECT  5.40 13.50 6.60 28.20 ;
        RECT  0.60 13.50 1.80 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.30 1.50 24.90 ;
        RECT  0.90 22.80 1.50 23.40 ;
        RECT  0.90 21.30 1.50 21.90 ;
        RECT  0.90 19.80 1.50 20.40 ;
        RECT  0.90 18.30 1.50 18.90 ;
        RECT  0.90 16.80 1.50 17.40 ;
        RECT  0.90 15.30 1.50 15.90 ;
        RECT  0.90 13.80 1.50 14.40 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 10.20 5.10 10.80 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 18.30 6.30 18.90 ;
        RECT  5.70 16.80 6.30 17.40 ;
        RECT  5.70 15.30 6.30 15.90 ;
        RECT  5.70 13.80 6.30 14.40 ;
        RECT  5.70 6.60 6.30 7.20 ;
        RECT  5.70 5.10 6.30 5.70 ;
        RECT  5.70 3.60 6.30 4.20 ;
        RECT  5.70 2.10 6.30 2.70 ;
        RECT  6.00 10.20 6.60 10.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 13.50 8.70 14.10 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 3.90 8.70 4.50 ;
        RECT  8.10 2.40 8.70 3.00 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.50 24.30 11.10 24.90 ;
        RECT  10.50 22.80 11.10 23.40 ;
        RECT  10.50 21.30 11.10 21.90 ;
        RECT  10.50 19.80 11.10 20.40 ;
        RECT  10.50 18.30 11.10 18.90 ;
        RECT  10.50 16.80 11.10 17.40 ;
        RECT  10.50 15.30 11.10 15.90 ;
        RECT  10.50 13.80 11.10 14.40 ;
        RECT  10.50 6.60 11.10 7.20 ;
        RECT  10.50 5.10 11.10 5.70 ;
        RECT  10.50 3.60 11.10 4.20 ;
        RECT  10.50 2.10 11.10 2.70 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.90 24.00 13.50 24.60 ;
        RECT  12.90 22.50 13.50 23.10 ;
        RECT  12.90 21.00 13.50 21.60 ;
        RECT  12.90 19.50 13.50 20.10 ;
        RECT  12.90 18.00 13.50 18.60 ;
        RECT  12.90 16.50 13.50 17.10 ;
        RECT  12.90 15.00 13.50 15.60 ;
        RECT  12.90 13.50 13.50 14.10 ;
        RECT  12.90 6.90 13.50 7.50 ;
        RECT  12.90 5.40 13.50 6.00 ;
        RECT  12.90 3.90 13.50 4.50 ;
        RECT  12.90 2.40 13.50 3.00 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  15.30 24.30 15.90 24.90 ;
        RECT  15.30 22.80 15.90 23.40 ;
        RECT  15.30 21.30 15.90 21.90 ;
        RECT  15.30 19.80 15.90 20.40 ;
        RECT  15.30 18.30 15.90 18.90 ;
        RECT  15.30 16.80 15.90 17.40 ;
        RECT  15.30 15.30 15.90 15.90 ;
        RECT  15.30 13.80 15.90 14.40 ;
        RECT  15.30 6.60 15.90 7.20 ;
        RECT  15.30 5.10 15.90 5.70 ;
        RECT  15.30 3.60 15.90 4.20 ;
        RECT  15.30 2.10 15.90 2.70 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        LAYER metal1 ;
        RECT  3.00 9.90 6.90 11.10 ;
        RECT  3.00 2.10 4.20 24.90 ;
    END
END BUFX8

MACRO BUFX4
    CLASS CORE ;
    FOREIGN BUFX4 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.00 10.80 3.60 11.40 ;
        LAYER metal2 ;
        RECT  2.70 10.50 4.20 11.70 ;
        RECT  3.00 9.90 4.20 11.70 ;
        LAYER metal1 ;
        RECT  2.70 10.50 3.90 11.70 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 5.40 6.30 6.00 ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 13.50 6.30 14.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 16.50 6.30 17.10 ;
        RECT  5.70 18.00 6.30 18.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 24.00 6.30 24.60 ;
        LAYER metal2 ;
        RECT  5.40 2.10 6.60 24.90 ;
        LAYER metal1 ;
        RECT  5.40 2.10 6.60 7.80 ;
        RECT  5.40 13.20 6.60 24.90 ;
        END
    END Y
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 10.80 1.20 ;
        RECT  7.80 -1.20 9.00 7.50 ;
        RECT  3.00 -1.20 4.20 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 10.80 28.20 ;
        RECT  7.80 13.50 9.00 28.20 ;
        RECT  3.00 13.50 4.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.00 10.80 3.60 11.40 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 16.80 3.90 17.40 ;
        RECT  3.30 15.30 3.90 15.90 ;
        RECT  3.30 13.80 3.90 14.40 ;
        RECT  3.30 6.60 3.90 7.20 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.40 9.00 6.00 9.60 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 18.00 6.30 18.60 ;
        RECT  5.70 16.50 6.30 17.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 5.40 6.30 6.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 9.00 7.50 9.60 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.30 8.70 24.90 ;
        RECT  8.10 22.80 8.70 23.40 ;
        RECT  8.10 21.30 8.70 21.90 ;
        RECT  8.10 19.80 8.70 20.40 ;
        RECT  8.10 18.30 8.70 18.90 ;
        RECT  8.10 16.80 8.70 17.40 ;
        RECT  8.10 15.30 8.70 15.90 ;
        RECT  8.10 13.80 8.70 14.40 ;
        RECT  8.10 6.60 8.70 7.20 ;
        RECT  8.10 5.10 8.70 5.70 ;
        RECT  8.10 3.60 8.70 4.20 ;
        RECT  8.10 2.10 8.70 2.70 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        LAYER metal1 ;
        RECT  0.60 8.70 7.80 9.60 ;
        RECT  5.10 8.70 7.80 9.90 ;
        RECT  0.60 2.10 1.80 24.90 ;
    END
END BUFX4

MACRO BUFX2
    CLASS CORE ;
    FOREIGN BUFX2 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 7.20 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.00 10.80 3.60 11.40 ;
        LAYER metal2 ;
        RECT  2.70 10.50 4.20 11.70 ;
        RECT  3.00 9.90 4.20 11.70 ;
        LAYER metal1 ;
        RECT  2.70 10.50 3.90 11.70 ;
        END
    END A
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 5.40 6.30 6.00 ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 13.50 6.30 14.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 16.50 6.30 17.10 ;
        RECT  5.70 18.00 6.30 18.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 24.00 6.30 24.60 ;
        LAYER metal2 ;
        RECT  5.40 2.10 6.60 24.90 ;
        LAYER metal1 ;
        RECT  5.40 2.10 6.60 7.80 ;
        RECT  5.40 13.20 6.60 24.90 ;
        END
    END Y
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 8.40 1.20 ;
        RECT  3.00 -1.20 4.20 7.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 8.40 28.20 ;
        RECT  3.00 13.50 4.20 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 3.90 1.50 4.50 ;
        RECT  0.90 2.40 1.50 3.00 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.00 10.80 3.60 11.40 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 18.30 3.90 18.90 ;
        RECT  3.30 16.80 3.90 17.40 ;
        RECT  3.30 15.30 3.90 15.90 ;
        RECT  3.30 13.80 3.90 14.40 ;
        RECT  3.30 6.60 3.90 7.20 ;
        RECT  3.30 5.10 3.90 5.70 ;
        RECT  3.30 3.60 3.90 4.20 ;
        RECT  3.30 2.10 3.90 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.40 10.50 6.00 11.10 ;
        RECT  5.40 9.00 6.00 9.60 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 18.00 6.30 18.60 ;
        RECT  5.70 16.50 6.30 17.10 ;
        RECT  5.70 15.00 6.30 15.60 ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 5.40 6.30 6.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        LAYER metal1 ;
        RECT  0.60 8.70 6.30 9.60 ;
        RECT  5.10 8.70 6.30 11.40 ;
        RECT  0.60 2.10 1.80 24.90 ;
    END
END BUFX2

MACRO AOI22X1
    CLASS CORE ;
    FOREIGN AOI22X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 12.00 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  8.10 5.40 8.70 6.00 ;
        RECT  8.10 6.90 8.70 7.50 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        LAYER metal2 ;
        RECT  7.80 5.10 9.00 21.90 ;
        LAYER metal1 ;
        RECT  5.40 5.10 9.00 7.80 ;
        RECT  5.40 2.10 6.60 7.80 ;
        RECT  7.80 19.20 9.00 24.90 ;
        END
    END Y
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  10.50 10.20 11.10 10.80 ;
        LAYER metal2 ;
        RECT  10.20 6.90 11.40 11.10 ;
        LAYER metal1 ;
        RECT  10.20 9.90 11.40 11.10 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 13.20 6.30 13.80 ;
        LAYER metal2 ;
        RECT  5.40 12.90 6.60 17.10 ;
        LAYER metal1 ;
        RECT  5.40 12.90 8.10 14.10 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 10.20 1.50 10.80 ;
        LAYER metal2 ;
        RECT  0.60 9.90 1.80 11.10 ;
        LAYER metal1 ;
        RECT  0.60 9.90 1.80 11.10 ;
        END
    END C
    PIN D
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 13.20 3.90 13.80 ;
        LAYER metal2 ;
        RECT  3.00 12.90 4.20 14.10 ;
        LAYER metal1 ;
        RECT  3.00 12.90 4.20 14.10 ;
        END
    END D
    PIN vdd!
        DIRECTION INPUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 13.20 28.20 ;
        RECT  3.00 19.50 4.20 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INPUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 13.20 1.20 ;
        RECT  10.20 -1.20 11.40 7.50 ;
        RECT  0.60 -1.20 1.80 7.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 10.20 1.50 10.80 ;
        RECT  0.90 6.60 1.50 7.20 ;
        RECT  0.90 5.10 1.50 5.70 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.30 3.90 24.90 ;
        RECT  3.30 22.80 3.90 23.40 ;
        RECT  3.30 21.30 3.90 21.90 ;
        RECT  3.30 19.80 3.90 20.40 ;
        RECT  3.30 13.20 3.90 13.80 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.00 6.30 24.60 ;
        RECT  5.70 22.50 6.30 23.10 ;
        RECT  5.70 21.00 6.30 21.60 ;
        RECT  5.70 19.50 6.30 20.10 ;
        RECT  5.70 6.90 6.30 7.50 ;
        RECT  5.70 5.40 6.30 6.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.20 13.20 7.80 13.80 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  10.50 24.00 11.10 24.60 ;
        RECT  10.50 22.50 11.10 23.10 ;
        RECT  10.50 21.00 11.10 21.60 ;
        RECT  10.50 19.50 11.10 20.10 ;
        RECT  10.50 10.20 11.10 10.80 ;
        RECT  10.50 6.60 11.10 7.20 ;
        RECT  10.50 5.10 11.10 5.70 ;
        RECT  10.50 3.60 11.10 4.20 ;
        RECT  10.50 2.10 11.10 2.70 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        LAYER metal1 ;
        RECT  0.60 17.40 11.40 18.30 ;
        RECT  0.60 17.40 1.80 24.90 ;
        RECT  5.40 17.40 6.60 24.90 ;
        RECT  10.20 17.40 11.40 24.90 ;
    END
END AOI22X1

MACRO AOI21X1
    CLASS CORE ;
    FOREIGN AOI21X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 9.60 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  5.70 2.40 6.30 3.00 ;
        RECT  5.70 3.90 6.30 4.50 ;
        RECT  5.70 5.40 6.30 6.00 ;
        LAYER metal2 ;
        RECT  5.40 2.10 6.60 6.30 ;
        LAYER metal1 ;
        RECT  3.00 2.10 6.60 6.30 ;
        RECT  0.60 8.10 4.20 9.00 ;
        RECT  3.00 2.10 4.20 9.00 ;
        RECT  0.60 8.10 1.80 24.90 ;
        END
    END Y
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  8.10 10.20 8.70 10.80 ;
        LAYER metal2 ;
        RECT  7.80 9.90 9.00 14.10 ;
        LAYER metal1 ;
        RECT  6.60 9.90 9.00 11.10 ;
        END
    END B
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 10.20 3.90 10.80 ;
        LAYER metal2 ;
        RECT  3.00 9.90 4.20 11.10 ;
        LAYER metal1 ;
        RECT  3.00 9.90 5.40 11.10 ;
        END
    END A
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  0.90 6.30 1.50 6.90 ;
        LAYER metal2 ;
        RECT  0.60 6.00 1.80 8.10 ;
        LAYER metal1 ;
        RECT  0.60 6.00 1.80 7.20 ;
        END
    END C
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 10.80 1.20 ;
        RECT  7.50 -1.20 8.70 7.50 ;
        RECT  0.60 -1.20 1.80 4.50 ;
        END
    END gnd!
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 10.80 28.20 ;
        RECT  5.40 15.00 6.60 28.20 ;
        END
    END vdd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  0.90 24.00 1.50 24.60 ;
        RECT  0.90 22.50 1.50 23.10 ;
        RECT  0.90 21.00 1.50 21.60 ;
        RECT  0.90 19.50 1.50 20.10 ;
        RECT  0.90 18.00 1.50 18.60 ;
        RECT  0.90 16.50 1.50 17.10 ;
        RECT  0.90 15.00 1.50 15.60 ;
        RECT  0.90 13.50 1.50 14.10 ;
        RECT  0.90 6.30 1.50 6.90 ;
        RECT  0.90 3.60 1.50 4.20 ;
        RECT  0.90 2.10 1.50 2.70 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 18.00 3.90 18.60 ;
        RECT  3.30 16.50 3.90 17.10 ;
        RECT  3.30 15.00 3.90 15.60 ;
        RECT  3.30 13.50 3.90 14.10 ;
        RECT  3.30 6.90 3.90 7.50 ;
        RECT  3.30 5.40 3.90 6.00 ;
        RECT  3.30 3.90 3.90 4.50 ;
        RECT  3.30 2.40 3.90 3.00 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 10.20 5.10 10.80 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 18.30 6.30 18.90 ;
        RECT  5.70 16.80 6.30 17.40 ;
        RECT  5.70 15.30 6.30 15.90 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 10.20 7.50 10.80 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  7.80 6.60 8.40 7.20 ;
        RECT  7.80 5.10 8.40 5.70 ;
        RECT  7.80 3.60 8.40 4.20 ;
        RECT  7.80 2.10 8.40 2.70 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  8.10 18.00 8.70 18.60 ;
        RECT  8.10 16.50 8.70 17.10 ;
        RECT  8.10 15.00 8.70 15.60 ;
        RECT  8.10 13.50 8.70 14.10 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        LAYER metal1 ;
        RECT  3.00 12.90 9.00 14.10 ;
        RECT  3.00 12.90 4.20 24.90 ;
        RECT  7.80 12.90 9.00 24.90 ;
    END
END AOI21X1

MACRO AND3X1
    CLASS CORE ;
    FOREIGN AND3X1 0 0 ;
    ORIGIN 0.00 0.00 ;
    SIZE 16.80 BY 27.00 ;
    SYMMETRY X Y ;
    SITE core ;
    PIN A
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  3.30 15.60 3.90 16.20 ;
        LAYER metal2 ;
        RECT  3.00 15.30 4.20 20.10 ;
        LAYER metal1 ;
        RECT  3.00 15.30 4.20 16.50 ;
        END
    END A
    PIN B
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  5.70 13.20 6.30 13.80 ;
        LAYER metal2 ;
        RECT  5.40 12.90 6.60 14.10 ;
        LAYER metal1 ;
        RECT  5.40 12.90 6.60 14.10 ;
        END
    END B
    PIN C
        DIRECTION INPUT ;
        PORT
        LAYER via ;
        RECT  10.50 16.20 11.10 16.80 ;
        LAYER metal2 ;
        RECT  10.20 15.90 11.40 17.10 ;
        LAYER metal1 ;
        RECT  10.20 15.90 11.40 17.10 ;
        END
    END C
    PIN Y
        DIRECTION OUTPUT ;
        PORT
        LAYER via ;
        RECT  15.30 7.20 15.90 7.80 ;
        LAYER metal2 ;
        RECT  15.00 6.90 16.20 8.10 ;
        LAYER metal1 ;
        RECT  14.10 6.90 16.20 8.10 ;
        RECT  14.10 2.10 15.30 24.90 ;
        END
    END Y
    PIN vdd!
        DIRECTION INOUT ;
        USE POWER ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 25.80 18.00 28.20 ;
        RECT  10.20 19.50 12.90 28.20 ;
        RECT  5.40 19.50 6.60 28.20 ;
        END
    END vdd!
    PIN gnd!
        DIRECTION INOUT ;
        USE GROUND ;
        SHAPE ABUTMENT ;
        PORT
        LAYER metal1 ;
        RECT  -1.20 -1.20 18.00 1.20 ;
        RECT  11.70 -1.20 12.90 4.50 ;
        RECT  3.90 -1.20 5.10 10.50 ;
        END
    END gnd!
    OBS
        LAYER cc ;
        RECT  -0.30 26.70 0.30 27.30 ;
        RECT  -0.30 -0.30 0.30 0.30 ;
        RECT  2.10 26.70 2.70 27.30 ;
        RECT  2.10 -0.30 2.70 0.30 ;
        RECT  3.30 24.00 3.90 24.60 ;
        RECT  3.30 22.50 3.90 23.10 ;
        RECT  3.30 21.00 3.90 21.60 ;
        RECT  3.30 19.50 3.90 20.10 ;
        RECT  3.30 15.60 3.90 16.20 ;
        RECT  4.20 9.60 4.80 10.20 ;
        RECT  4.20 8.10 4.80 8.70 ;
        RECT  4.20 6.60 4.80 7.20 ;
        RECT  4.20 5.10 4.80 5.70 ;
        RECT  4.20 3.60 4.80 4.20 ;
        RECT  4.20 2.10 4.80 2.70 ;
        RECT  4.50 26.70 5.10 27.30 ;
        RECT  4.50 -0.30 5.10 0.30 ;
        RECT  5.70 24.30 6.30 24.90 ;
        RECT  5.70 22.80 6.30 23.40 ;
        RECT  5.70 21.30 6.30 21.90 ;
        RECT  5.70 19.80 6.30 20.40 ;
        RECT  5.70 13.20 6.30 13.80 ;
        RECT  6.90 26.70 7.50 27.30 ;
        RECT  6.90 -0.30 7.50 0.30 ;
        RECT  8.10 24.00 8.70 24.60 ;
        RECT  8.10 22.50 8.70 23.10 ;
        RECT  8.10 21.00 8.70 21.60 ;
        RECT  8.10 19.50 8.70 20.10 ;
        RECT  9.30 26.70 9.90 27.30 ;
        RECT  9.30 -0.30 9.90 0.30 ;
        RECT  9.60 9.90 10.20 10.50 ;
        RECT  9.60 8.40 10.20 9.00 ;
        RECT  9.60 6.90 10.20 7.50 ;
        RECT  9.60 5.40 10.20 6.00 ;
        RECT  9.60 3.90 10.20 4.50 ;
        RECT  9.60 2.40 10.20 3.00 ;
        RECT  10.50 24.30 11.10 24.90 ;
        RECT  10.50 22.80 11.10 23.40 ;
        RECT  10.50 21.30 11.10 21.90 ;
        RECT  10.50 19.80 11.10 20.40 ;
        RECT  10.50 16.20 11.10 16.80 ;
        RECT  11.70 26.70 12.30 27.30 ;
        RECT  11.70 -0.30 12.30 0.30 ;
        RECT  12.00 24.30 12.60 24.90 ;
        RECT  12.00 22.80 12.60 23.40 ;
        RECT  12.00 21.30 12.60 21.90 ;
        RECT  12.00 19.80 12.60 20.40 ;
        RECT  12.00 10.20 12.60 10.80 ;
        RECT  12.00 3.60 12.60 4.20 ;
        RECT  12.00 2.10 12.60 2.70 ;
        RECT  14.10 26.70 14.70 27.30 ;
        RECT  14.10 -0.30 14.70 0.30 ;
        RECT  14.40 24.00 15.00 24.60 ;
        RECT  14.40 22.50 15.00 23.10 ;
        RECT  14.40 21.00 15.00 21.60 ;
        RECT  14.40 19.50 15.00 20.10 ;
        RECT  14.40 3.90 15.00 4.50 ;
        RECT  14.40 2.40 15.00 3.00 ;
        RECT  16.50 26.70 17.10 27.30 ;
        RECT  16.50 -0.30 17.10 0.30 ;
        LAYER metal1 ;
        RECT  9.30 2.10 10.50 11.10 ;
        RECT  7.80 9.90 12.90 11.10 ;
        RECT  3.00 17.40 9.00 18.60 ;
        RECT  3.00 17.40 4.20 24.90 ;
        RECT  7.80 9.90 9.00 24.90 ;
    END
END AND3X1

END LIBRARY
